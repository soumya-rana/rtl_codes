///////////////////////////////////////////////////////////////////////////////
// Company: Indian Institute of Science, Bengaluru 
// Engineer: Soumya Kanta Rana 
//
// Create Date: 17.11.2021
// Module Name: images ROM
// Project Name: ELM engine
// Target Devices: xc7a200tfbg484-2
//
////////////////////////////////////////////////////////////////////////////////
module test_images(input [8:0] addr,  output reg [255:0] data);
  always @ (addr) begin 
     case(addr)
      9'd1: data <=256'b0000000000111111000000001111000100000001110000000000001110000000000011110000000000011100000000000011100000000000011100000000000011110000000000001110011100000000111111111100000011100000110000001110000011000000111100001100000011111111100000000000010000000000; 
      9'd2: data <=256'b0111111111111100111000000000111100000000000001110000000111111110000000110000000000000011000000000000000111100000000000000111000000000000000110000000000000001110000000000000011100110000000000110011000000000011000110000000011000001111111111100000000111100000; 
      9'd3: data <=256'b0111111111000000111000001111000011000000001110001110000000011000011110000001100000011100011110000000111111111000000001111111000000011100111100000001110000111100000110000000110000011000000001100001110000000011000011100000001100000011110011110000000011111100; 
      9'd4: data <=256'b0000000001111111000000011110001100000111100000000000111000000000000111000000000000111000000000000111000000000000111000000000000011100000110000001100011111111100110011000001111011001100000001101110000000000110011100000001111000111111111111000000011111100000; 
      9'd5: data <=256'b0000111100000000000111100000000000111110000000000011111000000000001111100000000000111100000000000011111000000000001111100000000000011110000000000001111100000000000011110000000000001111100000000000011110000000000001111100000000000011111110000000001111110000; 
      9'd6: data <=256'b0000000000000110000000000000111000000000000011100000000000001100000000000000110000000000001111000000000011101100000000011100110000000111100111000001111000011000111110000000110011000000000110000000000000011000000000000000111100000000000011110000000000001110; 
      9'd7: data <=256'b0000011110000000000000011100000000000000111100000000000000110000000000000011100000000000001110000000000001100000000000001110000000000111110000000000111100000000011111000000000111110000000000111100000000000110110000000011111011110001111100000111111111000000; 
      9'd8: data <=256'b0000000000011000000000000111100000000000111100000000000111100000000000111000000000000111000000000001111000000000001110000000000001110000000001111110000000011110110000011111110011111111100111000000000000011000000000000011100000000000001110000000000000011100; 
      9'd9: data <=256'b0000111111111111001111100011111011111000001111101110000011111100111111111111110001111100001111000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000; 
      9'd10: data <=256'b0000100000000000000110000000000000011000000000000011100000000000001100000000000000110000000000000110000000000100011000000000111011000000001111111111111111111100111110000000110011000000000011000000000000011100000000000001100000000000000110000000000000011000; 
      9'd11: data <=256'b0000000000000001000000000000001100000000000001110000000000000110000000000000111000000000000111000000000000011100000000000011110000000000011110000000000011011000000000011001100000000111000100000000110000010000001110000001000011110000000000001000000000000000; 
      9'd12: data <=256'b0011111110000000111110111100000011110000111000000111111111100000001110001110000000000001110000000000001110000000000000111000000000000111000000000000111000000000000111000000000000111000000000000111000000000000111100000001111111111111111111000111111110000000; 
      9'd13: data <=256'b0001111111110000001100000001100001110000000011000110000000000110110000000000001111000000000000111100000000000011100000000000000110000000000000111000000000000011100000000000001011000000000001101110000000001100111100000011100000111001011000000001111111000000; 
      9'd14: data <=256'b1111111111100000110000000111000000000000001100000000000000110000000000000111000000000001110000000000011100000000000001110000000000000111111111000000000000011110000000000000011100000000000000110000000000000011000000000000011100000011111111100000001111110000; 
      9'd15: data <=256'b0000001111000000000001111000000000000110000000000001111000000000001110000000000001111000000000000111000000000000111000000000000011100000000000001110111111111100111011000000111011100000000001111111000000000111011110000000111000111111111111100000111111111000; 
      9'd16: data <=256'b0000111111111100000111000000111100111000000001110011100000000011001110000000011100111000000001110001110000001111000011100000110000000111111111000000111111111000111111001111000011000000001110001100000000011100111100000000110001111111111111000000111111111000; 
      9'd17: data <=256'b0000000000001110000000000001111000000000001110000000000001110000000000011110000000000011110000000000111100000000000111100000000000011100000000000111100000000000111100000001111011100000001111101111111111111110111111100001111000000000000011100000000000001111; 
      9'd18: data <=256'b0000000111111110001000000000011101110000000000110011100000111111001111111110000000011110000000000111111000000000111001100000000011000111100000001000000111000000110000001100000011100000111100000111100000111000000010000001100000001111111110000000000011110000; 
      9'd19: data <=256'b1110000001110000111110001111000001111111111100000111011111100000000000011000000000000011100000001100001100000000111111110000000001111111111111110011111000000000001111100000000000011110000000000000111000000000000011100000000000000110000000000000011000000000; 
      9'd20: data <=256'b0000000011110000000000011000000000000011000000000000011000000000000111000000000000011000000000000011000000000000011100011111110011101111100011111101100000000011111100000000001111100000000000111100000000000111011000000000111001111000011110000001111111100000; 
      9'd21: data <=256'b0000000000000111000000000000011100000000000011100000000000001110000000000000111000000000001111100000000000111110000000000111111000000001111011100000001110001110111111110000111000000000000011100000000000001110000000000000011000000000000001100000000000000010; 
      9'd22: data <=256'b0000111111111111001111000111111111110000000011111100000011111110111111111110111000000000000011000000000000011100000000000001100000000000001110000000000001111000000000000111000000000000111000000000000011100000000000001110000000000000111000000000000011000000; 
      9'd23: data <=256'b0000111111111100001110000000111001110000000001110110000000000111010000000000111000000000001111000001111111111000001111001111000001110000001110001100000000011100110000000000011011000000000001111110000000000011011110000000001100011111000001110000001111111100; 
      9'd24: data <=256'b0000011111111110001111100000011111111000000001111110000000000111110000000000111011000000001111101110000001111110011111111111110000111110011110000000000001110000000000001110000000000001110000000000001111000000000000111000000000000011100000000000001100000000; 
      9'd25: data <=256'b1111111111100000111000000111000000000000011100000000000001110000000000001110000000000001111000000001111111111100000011100000111000000000000001110000000000000011000000000000001100000000000000110000000000000011000110000000011100011111111111100000011111111000; 
      9'd26: data <=256'b0001111111111111000100000000000001110000000000001100000000000000110000000000000010000000000000001111000000000000011111100000000000000111100000000000000110000000000000011000000000000001100000000000000110000000000000111000000011111111000000000011110000000000; 
      9'd27: data <=256'b0000000111000000000011111111000000011110011110000011100000011100001100000000111001110000000001101110000000000111110000000000011111000000000001111100000000000110110000000000111011100000000111001111000001111000011111111110000000011111100000000000000000000000; 
      9'd28: data <=256'b0000111111100000000111111111000001111100011110001110000000111000110000000011100010000000001110000000000000111000000000000111000000000001111100000000011111000000011111111000000011111000000000001110000000000000111111111111111101111111111111100000011110000000; 
      9'd29: data <=256'b0000001111111111000000000000000000001110000000000001110000000000011110000000000011100000000000001111111111110000000000000111100000000000000111000000000000001110000000000000111000000000000111000111000000111100011000000111000001111111111000000001111100000000; 
      9'd30: data <=256'b1111111000000000000011111100000000000000111000000000000011100000000000001100000000000001110000000000011111111111000111111111111000111111100000000000011100000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000; 
      9'd31: data <=256'b0001111111111000011111000000000011000000000000001100000000000000111000000000000001111000000000000001110000000000000011111100000000000001111110000000000000011100000000000000111100000000000000110000000000000011010000000000001101111111111111110000000111111000; 
      9'd32: data <=256'b0001111111111100000000000000110000000000000011100000000000001100000000000001110000000000001110000000000001110000000000001100000000011111111111100001111111111111000111110001000000011100000000000111100000000000011100000000000011110000000000001100000000000000; 
      9'd33: data <=256'b0000000000111111111111111111111001111111111100000000000111000000000001111000000000001111000000000011110000000000001111111110000000111111111111000000000000011110000000000000011000000000000011100000000000011100000000001111100001111111111000000111110000000000; 
      9'd34: data <=256'b0000111111000000000111111111110001111000000011100111000000001110010000000000011100000000000000110000000000000011000000000000011100000000000001101100000000001110110000000001110011000000011110001111000111110000011111111100000000011110000000000000000000000000; 
      9'd35: data <=256'b0000000011111100000110000000001100110000000000110011000000000011000110000001111000011100001110000000111111110000000001111000000000000001110000000001100001110000111100000011100011000000000011001100000000001110111000000000011001111111111111100000001111111000; 
      9'd36: data <=256'b0000011111111000000111111011110000111110000001100111000000000011011100000000001101100000000000110111110000000011011110000000011101110000000001100111000000001110111110000001110011111111011110001100000111110000111111111100000001111111000000000011110000000000; 
      9'd37: data <=256'b0000111000000000001110000000000111100000000000111100000000001110110000000111110011101111111000001111111111111111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000111000000000000011100000000000000110; 
      9'd38: data <=256'b0000011111111111000001111111000011100000000000001100000000000000110000000000000011000000000000001110000000000000001100000000000000011110000000000000001110000000000000011100000000000000011000000000000011100000000000001100000000111111100000000000111000000000; 
      9'd39: data <=256'b0011111111111100011110000000111011100000000001101100000000001110111110000111110001111111111111100011111111111111000000000000011100000000000001110000000000000111000000000000011100000000000001100000000000001110000000000001111000000000000011100000000000000100; 
      9'd40: data <=256'b0000000011111111000011111110000000011110000000000011110000000000001110000000000000110000000000000011000000000000001111111110000000111100011111100000000000000011000000000000001100000000000000110000000000001110000000000000110011000001111110001111111110000000; 
      9'd41: data <=256'b0000000011100000000000001110000000000001111000000000001111100000000000111111000000000111111100000000011101110000000011100011100000111100001111000111000000011100111000000001110011100000000011100000000000000110000000000000011000000000000000100000000000000011; 
      9'd42: data <=256'b1000000000111000111111111111100000001111111000000000000011100000000000001100000000000000110000000000000111000000000000011000001000011111111111110000111110000000000000011000000000000001100000000000000110000000000000011000000000000000110000000000000010000000; 
      9'd43: data <=256'b0000111011100000000111001111000000111000011111110110000000001111111000000000000011000000000000001110000000000000111000000000000011111110000000000001111110000000000000111000000000000011100000000000001110000000010111110000000001111000000000000011000000000000; 
      9'd44: data <=256'b0001111111111100001111111000111011111000000001101111100000000111111100000000011111110000000001101111000000000110111000000000111011100000000111101110000000011100111000000011100001110000011100000111000011100000011111111100000000111111100000000000011000000000; 
      9'd45: data <=256'b0000111111000000000110001110000000000000111000000000000111000000000001111000000000001111111100000000000000111100000000000000111100001111000000110000000000000011000000000000001111000000000000111110000000000110011111000000111000001111111111000000000111110000; 
      9'd46: data <=256'b0000011100000000000001110000000000000110000000000000111000000000000011000000000000011100000000000011100000000000011100000000000011100000000011111100000000001111110000000000111111000000001111101111111111111110000111000000111000000000000001100000000000000111; 
      9'd47: data <=256'b0000011111111000000011111111100000000000001110000000000001110000000000001111000000000111111111000000011111111110000000000000111100000000000001110000000000000111000000000000011100000000000011110111111000011110111100011111110011111111111100001111111110000000; 
      9'd48: data <=256'b0001111111111100000000000000111000000000000001110000000000001110000000001111110000000011111000000000111100000000000001111000000000000001111100000000000000110000000000000011100000000000001110001110000001110000111000011110000001111111110000000001110000000000; 
      9'd49: data <=256'b0001100000000000000110000000000000011000000000000001100000000000001100000000001100110000000001110111000000000111011000000000011101100000000001101100000000000110110000011111111011111111110111100000000000000110000000000000011000000000000011000000000000001100; 
      9'd50: data <=256'b0111111110000000110000011111000000000000001110000000000000011000000000000001100000001111111110000001111111111000000011110111111000000000000001110000000000000011000000000000001100000000000000111110000000000111111100000000111000111111111111000000001111100000; 
      9'd51: data <=256'b0000000001111110000000011100111100000011000011110000011000011111000001100011011000000011111011100000000000001100000000000011100000000000111100000000000111000000111111110000000011111100000000110000111000000111000001110000011000000011111111000000000001100000; 
      9'd52: data <=256'b0000000000011110000000000111100011111111111100000000000011100000000000001100000000000001100000000000001110000000000000110000000001111111110000001111111111111110100011100000111100001100000000000000110000000000000111000000000000011000000000000001100000000000; 
      9'd53: data <=256'b0001100000000000001110000000000001110000000000001111000000000000111000000000000011000000000000001100001111100000110111111111100011111111011111101110000000001111111000000000011111110000000001111111111000000111000111110000011100000111111111110000000000110000; 
      9'd54: data <=256'b0000011111110000000011100001000000111000000100000010000000000000001000000011111001100000111000100111111110000011001111000000001100000000000000110000000000000011000000000000001100000000000001100000000000000110111111000011110000011111111100000000000011000000; 
      9'd55: data <=256'b0000000000000001000000000000001100000000000001100000000000000110000000000000111000000000000111000000000000111000000000000111100000000001110110000000000110010000000001110011000000011100001000000111000000100000111000000110000000000000010000000000000011000000; 
      9'd56: data <=256'b0011111111110000011100000011100011000000000110000000000001111000000000001111000000000000111000000000001110000000000000111000000000000001111110000000000001111110000000000000001100000000000000110000000000000111000000000001110000010001111110000011111111000000; 
      9'd57: data <=256'b0000001111110000000011111111110000001100000011100001100000000110001110000000001111110000000000111110000000000011111000000000001111100000000000111111000000000011111110000000011001110000000011100011110000111100000111111111100000000111111000000000000000000000; 
      9'd58: data <=256'b0000000011111100000000000000110000000110000001100001110000000110001110000000011001110000000001110110000000000111111000000000011111100000000001111100000000000111111000000000111111100000000011101110000000011100011110000011110000111111111110000000111111100000; 
      9'd59: data <=256'b0000000000111111000000011111000000000111100000000000111000000000000111100000000000111000000000000111000000000000011000000000000011100011111100001100011000011100110000000000110011000000000011001110000000001100111100000001110000111111111110000000001111000000; 
      9'd60: data <=256'b0000011111111111001111110000000011111000000000001110000000000000111000000000000011110000000000000011111000000000000001111100000000000000011110000000000000001100000000000000011100000000000000110000000000001110000000000011110011111111111000000000111000000000; 
      9'd61: data <=256'b1100000000000000011100000011100001110000011111000001111111111000000011111111000000000011110000000000001100000000001111110000000000111111000000000000111111111100000011111111111100001100000000000000110000000000000111000000000000011100000000000001100000000000; 
      9'd62: data <=256'b0000000000001111000000000011100000000001111100000000001110000000000011110000000000111100000000000111000000000000011100000000000011100111111000001100110001100000111110000011000011110000011000001110000001100000111110011100000001111111000000000011111000000000; 
      9'd63: data <=256'b0011111111111100011101111111111101000000000000000000000000000000011000000000000011100000000000001100000000000000111000000000000011111000000000000011110000000000000011110000000000000011100000000000001110000000000001111000000011111110000000000011100000000000; 
      9'd64: data <=256'b0000000000000111000000000000011100000000000001110000000000000110000000000000011000000000000011100000000000001110000000000000111000000001100011000000001100001100000011100000110000111000000111000111000000011000110000000001100000000000000110000000000000011000; 
      9'd65: data <=256'b0111111111111111111111111000011111000000000011110100000000001110000000000011110000000000011110000000000011100000000000011111000001111111111110000111101110000000000001110000000000000111000000000000111000000000000001110000000000000111111100000000000011000000; 
      9'd66: data <=256'b0000011111111000000111100000111101111000000011110110000000011111011111111100111100011111000011101100000000001110110000000011111011000000111111101111111110000110001111000000011100000000000001110000000000000011000000000000011111111111111111100111000000000000; 
      9'd67: data <=256'b0000000111111111001111111111110001100000000000000000000000000000000000000000000000101111100000000111110111100000011100000110000001100000011000000110000001110000000000000011000000000000001100000000000001110000110000000110000001111110111000000000111111000000; 
      9'd68: data <=256'b0000000011111110000000011100011000000011100000110000000111000110000000000000111000000000000111000000000001110000000000011110000000011111100000001111110000000000001111100000000000001111100000000000000111000000000000001111000000000000001111000000000000001111; 
      9'd69: data <=256'b0000000001111110000000011111110000000011110000000000111110000000001111100000000000111000000000000111100000000000111100000000000011100000000000001110000000000000111000000000000011111111111111111111111000000111111111000000011101111111111111100000001111110000; 
      9'd70: data <=256'b0000000000000111011111111111111100001111110011100000000000011100000000000011100000000000011000000000000011100000000000001100000000111111111111111111111100000000000011100000000000011100000000000011100000000000001110000000000001111000000000000010000000000000; 
      9'd71: data <=256'b0000001111111110000000111000011100000011000000110000001100000110000000111001111000000001111110000000111011100000000001111000000000000111100000000000110011000000001110001110000001100000011000001100000011100000110000111100000011111110000000000110000000000000; 
      9'd72: data <=256'b0000011111111111111111111111111101111111000111110110000000011110011000000011110001111111111110000011111110111000000000000011000000000000001100000000000001110000000000000110000000000000111000000000000011100000000000001110000000000000111000000000000011000000; 
      9'd73: data <=256'b0000000000000111000000000001111100000000001111110000000011111110000000011110110000000111100111000000111100111000000111000011000001111100001100001111000001100000110000001110000000000000111000000000000011000000000000011000000000000000110000000000000011000000; 
      9'd74: data <=256'b0000000011111000000111111111000011111110000000001000000000000000110000000000000011110000000000000011111100000000000000111100000000000000111110000000000000011110000000000000011100000000000000110000000000000011011100000000111001111111111111000000111111000000; 
      9'd75: data <=256'b1111111100000000000011111000000000000001110000000000000011100000000000001110000011100001111000001111111111000000000111111110000000000000111110000000000000011110000000000000011000000000000001110000000000000111001110000000111100111111111111110000001111110000; 
      9'd76: data <=256'b0000011111111100000011110000011000011100000000110011100000000010000111000000011000011100000001100000111100011100011111111111100011100111111100001100111111110000110000000011111011000000000011111110000000000111011110000000011100011111000111100000001111111110; 
      9'd77: data <=256'b0011111100000000000000111000000000000001100000000000000110000000000000011000000000000011100000000000011100000000001111111000000000000000111100000000000000111000000000000000111000000000000000100000000000000011110000000000001111111110111111110000011001100000; 
      9'd78: data <=256'b0000000000111100000000001111100000000001111000000000011110000000000011110000000000011100000000000011110000000000011110000000000011100000011110001110011111111110110011110000011011111110000001111111000000000111111100000001111101111111111111000000011111100000; 
      9'd79: data <=256'b0000111111111111011110000000000101000000000000000100000000000000010000000000000011000000000000001111111100000000111111111110000000000000011110000000000000011000000000000000110000000000000001100000000000001100000000000001110000000011111110000000000110000000; 
      9'd80: data <=256'b0000011111111100000111110000111000011100000001100111100000000111011000000000001111101000000000111101100000000011110110000000001111011000000001111111100000000110011110000000111000111000000011000001110000111100000111000111100000001111111100000000011111000000; 
      9'd81: data <=256'b0000011110000000000111111000000000111111000000000111000000000000011100000000000011100000000000001110000000011100111000000011110011110000001111100111111111111110000001110000111000000000000011110000000000001111000000000000011100000000000000110000000000000011; 
      9'd82: data <=256'b1111111111111000000011110001100000000000001110000000000000110000000000000111000000000011110000000000011110000000001111111111000000111000001111000000000000001100000000000000111000000000000001110000000000000011000000000000001101111111111111110000001111111110; 
      9'd83: data <=256'b0000111111111100001111110000111001111100000011110111000000000111111000000000001111100000000000111100000000000011110000000000001111000000000001111100000000000110111000000000111011100000000111100111000000111100011111111111100000011111111000000000011110000000; 
      9'd84: data <=256'b1111111111110000110000000011100000000000000110000000000000011000000000000011000000001111111000000000001111000000000000001111110000000000000001110000000000000011000000000000011100000000000011000000000000011000011000001111000011111111100000001111110000000000; 
      9'd85: data <=256'b0000000000111110000000000111110000000000111100000000001111100000000001111000000000011111000000000001110000000000011110000000000001110000000000111110000000001111111000001111111011111111111111100111111100011110000000000001111000000000000111100000000000011111; 
      9'd86: data <=256'b0000000011111110000000111110111100001111100001110001111000000111011110000000011111110000000001111111000000000111111100000000111011100000000011100110000000011100011000000001110001100000001110000111000001110000011100011110000000111111110000000000111100000000; 
      9'd87: data <=256'b0000000011111111000000011100001100000011110000110000011110001110000011110001110000000111111110000000001110000000000001100000000000000110000000000000111000000000000011000000000000011000000000000011000000000000011000000000000011100000000000001100000000000000; 
      9'd88: data <=256'b0000000000000111000000000000111000000000000111100000000000111100000000001111110000000001100111000000011100011000000011000001100011111000000110001000000000110000000000000011000000000000011100000000000001110000000000001110000000000000111000000000000011000000; 
      9'd89: data <=256'b0000000000110000000000001110000000000001111000000000001110000000000001110000000000001110000000000011111000000000001110000000000011110000000011111111111111111111000111110011100000000000001110000000000001111000000000001111000000000000111110000000000001110000; 
      9'd90: data <=256'b1111111110000000100001111000000000000011100000000000000110000000000000111000000000111111100000000001101111100000000000001111000000000000001111000000000000001110000000000000111000000000000011110000000000001110000000000111110001111111111110001111111111000000; 
      9'd91: data <=256'b0000000001111000000000011110000000000011100000000000111100000000000111100000000000111000000000000111000000000000111000000000000011100000001111111100001111111110111111111011110001111110011110000000000011110000000000001100000000000001110000000000000011000000; 
      9'd92: data <=256'b0000111111111110000000000011000000000000000000000001110000000000000111111000000000011111111100000001110001111110000111000000011100000000000001110000000000000011000000000000001100000000000001111100000000011111111000000111110011111111111100000011111111000000; 
      9'd93: data <=256'b0000000011110000000000011100000000000111100000000000111000000000000111000000000000111000001100000111000000110000111000000011100011000000000111001100000000011100111111111111111000000000000001100000000000000111000000000000001100000000000000110000000000000011; 
      9'd94: data <=256'b0000000000111110000000111111111000000111000011000011110001111000000000011110000000000011000000000001111000000000011110000000000001111111111111100000000000001111000000000000001100000000000001110000000000001110111110000011110011110001111110001100001110000000; 
      9'd95: data <=256'b0000000011111111000111111111111111111000000111000000000000111000000000000111000000000000111000000000000011100000000000011000000000000011100000001111111111111111000011100000000000001110000000000001110000000000000110000000000000111000000000000011100000000000; 
      9'd96: data <=256'b0011111111111110111101110011111111011100000110111001100000011111111110000001111000111000001111000001111111111000000000000001100000000000001100000000000000110000000000000110000000000000011000000000000011100000000000001100000000000000110000000000000011000000; 
      9'd97: data <=256'b0000111111111100001111100001111001111000000011100110000000000011011000000000001111000000000000111100000000000011110000000000001111000000000001111100000000000110110000000001110011000000001111001110000000111000011100001111000000111111111000000001111110000000; 
      9'd98: data <=256'b0000011111110000001111110011100011100000000110000000000000111000000000000011000000000000001100000000000000110000000000000111011100011111111111110011111001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001000000; 
      9'd99: data <=256'b0111111111111100000000000001110000000000001110000000000001111000000000001111000000000000111000001111000111000000111110111000000000111111100000000001111111111100000111100011111100011100000000000001110000000000001110000000000000111000000000000011100000000000; 
      9'd100: data <=256'b1110000000111110011111111111110000011111111000000000000011000000000000011100000000000011100000000001111100000000001111111111111100001111111111110000011000000000000011100000000000001100000000000000110000000000000111000000000000011100000000000001111000000000; 
      9'd101: data <=256'b0000000000001110000000000001111000000000001111110000000001111110000000001111110000000001111111000000000110111100000001111011100000001111001111000001110000111101011110000011111111111000111111101111111111111100000000000001110000000000000111000000000000001100; 
      9'd102: data <=256'b0000000000111111000000011110000000000011100000000000011100000000000011100000000000011100000000000011100000000000001100000000000001110111111111101111111000000110111110000000011111110000000001101111000000001110111100000011110011111111111100000111111111100000; 
      9'd103: data <=256'b0000011111111100001111110000011001111000000001111111000000011111110000000001111011000000011111001111111111111100000011111111100000000000001110000000000000111000000000000011100000000000011100000000000011100000000000011100000000001111110000000000110000000000; 
      9'd104: data <=256'b0000000001111111000000001110000000000011110000000000111100000000000111100000000000111100000000000111100000000000111100000000000011100000000000001110001111111000111111111111111011101000000011101110000000001110111110000011111000111111111110000000111111000000; 
      9'd105: data <=256'b0000000111111111000111111100111011111100000111100000000000011000000000000111100000000000011100000000000011100000000011001100000000001111110000000000011111111111000000110011110000000111000000000000011000000000000011100000000000001110000000000000011000000000; 
      9'd106: data <=256'b0000000011111000000000111110000000000111110000000000111000000000001111100000000000111000000000000111000000000000011100000000000011100000000000001110011111110000111111111111110011111100000011101111100000001111011111100011111000111111111110000000001110000000; 
      9'd107: data <=256'b0000000011111111000000111100001100001111111001110000110000000110000011100001110000011110001110000000111101100000000001111110000000000111100000000000111111000000001111011110000001110000111000000110000011100000110000001110000011111111110000000011111000000000; 
      9'd108: data <=256'b0000001111111111000111100000011101111100000001110111000000001111111000000011111011100000011111000111111111101100001111110000110000000000000011000000000000001100000000000001110000000000000111000000000000111000100000000011100011111000011100000001111111100000; 
      9'd109: data <=256'b0000011111111110000001100111111000000000011110000000000011110000000000111110000000000111111100000000011111111110000001111111111000000000000011110000000000000111000000000000011100000000000001111100000000011110111111111111110011111111111110000011111110000000; 
      9'd110: data <=256'b0000000001111000000000001111000000000011111000000000011111000000000011111000000000011110000000000011110000000000011110000000011101111000000011101110000000011110111111111111111000000000001111000000000000111100000000000011100000000000001111000000000000001110; 
      9'd111: data <=256'b0000000011000000000000011110000000000011111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000001111000000000000111100000000000011110000000000011110000000000011111100000000000011111100000000000111000000; 
      9'd112: data <=256'b1111111111100000000000001111100000000000001110000000000000111100000000000011100000000000011100000011110001110000001111111111100000000011111111110000000111000000000000011000000000000011100000000000011100000000000001110000000000000111000000000000011100000000; 
      9'd113: data <=256'b0000001110000000000001110000000000001111000000000000110000000000000111000000000000011100000000000011100000000000001110000000000000111000100000000011111111111100001111000001111111111000000001111111110000000111000111000000111100001111111111100000000111110000; 
      9'd114: data <=256'b0000000000111111000000001111100000000011110000000000011100000000000011100000000000111100000000000011000000000000011100000000000011100000000000001100000000000000111111111111000011111100001111001100000000001100111100000001110001111111111110000000011110000000; 
      9'd115: data <=256'b0000111111111100000111000000110000111100000001100011100000000110111100000000011111100000000000111110000000000011110000000000001111000000000000111100000000000011110000000000011111000000000001111110000000001110011110000001110000111111111110000000011111000000; 
      9'd116: data <=256'b0111111111110000111100000111100000000000000110000000000000011100000000000001110000000000000110000000000000011000000000000011100000000000001110000111111111111111000000000111000000000000011000000000000011100000000000011100000000000111100000000000011000000000; 
      9'd117: data <=256'b0111111100000000111000011100000000000000110000000000000001100000000000001110000000000001110000000000001110000000011111110000000000000001111100000000000000111000000000000000111000000000000001101110000000000011011100000000001100111111110111100000011111111100; 
      9'd118: data <=256'b0000111111100000000111000001100000111000000011100110000000000110111000000000001111000000000000111100000000000011100000000000000110000000000000011000000000000011100000000000001111000000000001101100000000001100011000000011110000111000111100000001111111000000; 
      9'd119: data <=256'b0000111111100000111111101110000000000000110000000000000011000000000000001000000000000001100000000111001110000000111111111111100000000111011111110000111000000000000011000000000000001100000000000111110000000000011110000000000000111000000000000011100000000000; 
      9'd120: data <=256'b0011111111111100001110111111111100111000000000000011000000000000011000000000000001110000000000000011000000000000001111000000000000001111000000000000001111100000000000001110000000000000011100000000000001100000111110111110000011111111100000000001000000000000; 
      9'd121: data <=256'b0000001110000000000001110000000000011110000000000001110000000000011110000000001111100000000001111100000000001110110000000001111111111111111111000000000000111000000000000011100000000000011100000000000001110000000000000111000000000000011100000000000000110000; 
      9'd122: data <=256'b1111110000000000100011100000000000000111100000000000001110000000000000111100000000000011110000000000011110000000001111111111110000011000000111100000000000000111000000000000011100000000000011100000000000011110000000000111110000000011111100000000111111000000; 
      9'd123: data <=256'b0000000000111111000000001111110000000011100000000000111100000000000111000000000000111000000000000111000000000000111000000000000011100000000000001110000111100000110000110011000011000000001100001100000000110000111000000110000011111111111000000011111100000000; 
      9'd124: data <=256'b0000000000011100000000000111110000000001111100000000011111000000000011111000000000111110000000000111100000000000011111111111000001111111111111101111110000001111111110000000001111111000000000110111110000000111000111100000111100001111111111100000001111110000; 
      9'd125: data <=256'b0011111111110000011110000111100011110000000111001110000000001100111000000000111011000000000001111100000000000011110000000000001111000000000000111100000000000011111000000000001101110000000001110011100000001110001111000001111000001111111110000000011111110000; 
      9'd126: data <=256'b0001111111110000111111111110000011110001111000000000000111000000000000111000000000000111100000000000011110000000000001110000000000001111011111110111111111111100001111100000000000111100000000000111000000000000011100000000000011110000000000000110000000000000; 
      9'd127: data <=256'b0000000000011111000000001111000000000000111000000000001110000000000001110000000000001110000000000001110000000000001100000000000001110000011111101110000111100110110000110000011011001111000011101111110000111100111110000111000001111111111000000000010000000000; 
      9'd128: data <=256'b0011111111100000000000001111110000000000000111110000000000000111000000000001111000000000111111000000001111100000000000111100000000000001111110000000000000111110000000000000011100000000000111100000000011111100000001111110000000111111000000001111100000000000; 
      9'd129: data <=256'b0000111111111110000011000000011100111111100001110111000111100000111000001111111011111111111001110111110000000111000000000001110000000000001111000000000011111000000000011110000000000001110000000000001110000000000001110000000000000111110000000000000011110000; 
      9'd130: data <=256'b0000111111100000000111000111000000010110001110000011011000111000001111100011100000011110001110000000000000110000000000000111000000000000111100000000000011100000000000111100000000111111100000110110111100000011111111111100011111000000111111100000000000111000; 
      9'd131: data <=256'b0000000000000111000000000000111100000000000111100000000000011100000000000011100000000000111110000000001111110000000011100011000000111100001100001110000000110000000000000110000000000000011000000000000001100000000000000110000000000000001100000000000000011000; 
      9'd132: data <=256'b0000000000000011000000000000001100000000000001110000000000001110000000000000111000000000001111100000000000111100000000000110110000000001110011000000001110001100000011100000110000001100000011000001100000001100111100000000110011000000000011000000000000001110; 
      9'd133: data <=256'b0111111111110000000000111111110000000000000000001000000000000000100000000000000010000000000000001111100000001100000000000000011000000000000000110000000000000011000000000000001100000000000000110000000000000111000000000001110000011100011110000000111111110000; 
      9'd134: data <=256'b1100000000000111111100000001111000111111111110000000000000110000000000000111000000000000011000000000000011100000001111101100000000111111111111110001100011000000000010011100000000000001100000000000000110000000000000111000000000000011100000000000001110000000; 
      9'd135: data <=256'b0000000111110000000000111111000000001111101100000000111001100000000111100111000000011000000000000111100000000000011100000000000011110000000000001111111111111000111111100001111011110000000001101111100000000111011100000000111001111111111111100001111111100000; 
      9'd136: data <=256'b0001111111111110000010000000000000011000000000000001100000000000001100000000000000111111111110000011110000011110000100000000111000000000000000110000000000000011000000000000001100000000000000110000000000001110000000001111110011111111110000001111000000000000; 
      9'd137: data <=256'b0000011111111100000011111111000000011110011110000011111111111110001111110001110000111111001111000011111000111000001111111111100000001111111100000000001111100000000000001111100000000000001111000000000000011110000000000000011111111111111111111111000000011110; 
      9'd138: data <=256'b0111111111111000111000000000000011000000000000001100000000000000111000000000000001111110000000000000111100000000000000111100000000000000111110000000000001111000000000000001111100000000000001111100000000000011111100000000011111111111111111110000111111111110; 
      9'd139: data <=256'b0000011111100000000111110111100001111101101110001111111100011000110000111111100011100000111110001111111111111110001111111000111000000000000001110000000000000111000000000000011100000000000011110000000001111100000000111111100000111111110000000111110000000000; 
      9'd140: data <=256'b0000000111111100000111110011111000111000001110101110000000111011110000000011101110000000001110111100000000111110011000000111100001111111111110000000000000111000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000; 
      9'd141: data <=256'b0000111111111000001111100001111001111000000001110110000000000011011110000000011101111110000001101110001111111110111111111111110000111111110111000000000000011100000000000001110000000000000111000000000000011100000000000000110000000000000011000000000000001100; 
      9'd142: data <=256'b0001111111110000001110000011100001110000000010001110000000001100110000000000011010000000000001111000000000000011100000000000001110000000000000110000000000000011000000000000011000110000000001100011100000001110000111000001110000001111111110000000001111110000; 
      9'd143: data <=256'b0000000111000000000000111000000000000111100000000000111000000000000011100000000000111100000000000111100000000000011100000000000001100000000000101110000000001111111000011111111011111111000111000111100000011000000000000011100000000000000110000000000000011100; 
      9'd144: data <=256'b0000011110111000000011100000111000011110000001100011111000000111001110000000001101111000000000110111000000000011011100000000011111100000000001111100000000001110110000000011110011000000011110001100000111100000111001111100000011111111000000000011100000000000; 
      9'd145: data <=256'b0000000011000000000000111100000000001111110000000001110011000000011100001100000011100000110000001100000011000000100000001100000011100000110000110111111111111111000001111111100000000000100000000000000010000000000000001000000000000000100000000000000110000000; 
      9'd146: data <=256'b0000000001111000000000001111000000000000111000000000000111100000000000111100000000000111100000000000111100000000000011100011100000011111111111100011111111011110011111000011110011111100011110001111111111100111111111111111111011111111111110001111000000000000; 
      9'd147: data <=256'b0000000011111110000000001100011100011100000011100001100000011000000111100111100000000110111000000000001111000000000001111100000000001110111000000001110001110000001110000001100001110000000110001110000000011000011100001111100000111111110000000000010000000000; 
      9'd148: data <=256'b0111111111000000111000001110000000000000111000000000000011100000000000001100000000000011100000000001111110000000011111111110000001100000011111000000000000001110000000000000011100000000000001110000000000000111000000000000111111111111111111101111111111100000; 
      9'd149: data <=256'b0000000001110000000000111100000000000111100000000000111000000000000110000000000000110000000001110111000000000111111000000001111011100000001111001110000111111100111111111111100001111100001110000000000000111000000000000011100000000000011100000000000000110000; 
      9'd150: data <=256'b0000111111110000001111000011100001110000000010000110000000011000001110000011100000011100001100000000111101110000000000111100000000001111011100000111110000011100111000000000011011000000000001111000000000000011111000000000001100111111111111110000001111111000; 
      9'd151: data <=256'b0001111111111000001111000001111000110000000000110011100000000011000111000000011100001111000011110000011110111100111111111111100011111111110000001110000011100000011000001110000001100000011000000011000001100000000110000110000000011111111000000000011111000000; 
      9'd152: data <=256'b0000000111111111000000111100001100001111000000110001111000000011001110000000001100110000000000110110000000000011111000000000001011000000000000111100000000000011110000000000001111000000000011101100000000011110111100000111110001111111111100000001111111000000; 
      9'd153: data <=256'b0111111110000000011000111111000000000000011110000000000000011100000000000001110000000000001111000000000001111000000000001110000000000001111000000000011110000000000111100000000001111000000000001110000000000000110000000001111111111111111111100001110000000000; 
      9'd154: data <=256'b0000000111111110000000000000011100000000000001100011000000011110001100000011100000111000011100000001111111100000000001111100000000001111111000000011110001111000011100000001100011100000000110001110000000111000111000001111000011111111111000000111111111000000; 
      9'd155: data <=256'b0001111111100000001110001111000000110000001100000011111110111000000110111011100000001111001110000000000000110000000000000111011000000000111001110000000111000111000000111000001111001111000000111111110000000011001111111100001100000011111111110000000000111110; 
      9'd156: data <=256'b0000000000000111000000000000011100000000000001110000000000001110000000000000111000000000000111100000000001111110000000001111111000000001111011100000001110001100000011110000110000111100000111001111100000011100000000000001100000000000000110000000000000011000; 
      9'd157: data <=256'b0000001111111111000011110000001101111100000000110110000000000011110000000000011010000000000011000000000000111000000000000111000000000000110000000000011110000000000011100000000011111000000000001100000000000000111110000000110000011111111111000000011111110000; 
      9'd158: data <=256'b0001111111111100011100000000011001100000000000110110000000000011011100000000001100110000000001110001111000011110000001100111100000011111111000001111111111100000110000000011000011000000001110001110000000011000001110000001100000011111111110000000011111100000; 
      9'd159: data <=256'b0000011111110000000011000011100000011000111110000011000001111000001100000011100011111111111110001111111110011100000000000000111000000000000011100000000000000111000000000000001100000000000000110000000000000011000000000000111000000000011111000111111111110000; 
      9'd160: data <=256'b0000111111111100001111100001111001111000000011101111100000011110111000001111110011111111111111101111111111111110011111111000111000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111100000000000011110000000000001111; 
      9'd161: data <=256'b0000000000001111100001111111111011111111111111000000010001110000000000001110000000000000111000001111111111000000111111111111110001100111111111000010111100000000000011100000000000001110000000000001111000000000000111000000000000011100000000000001110000000000; 
      9'd162: data <=256'b0000000000111111000000000110000000000011110000000000001000000000000111100000000000011000000000000011000000000000011000000000000001100011111000001110111111111110110111000000011111111000000000111111000000000011111110000000011100111111111111000000111111110000; 
      9'd163: data <=256'b0000000001111000000000011111000000000111100000000000111000000000000111000000000000111000000000000111000000000000111000000001100011100011111111111100011100000111110001100000011111000000000001111100000000001110111000000011110001111111111100000000111100000000; 
      9'd164: data <=256'b0000011111111110000001100000001100000100000000010000011000000011000001110000011100000011100111000000000111111110000000111111100000011111111000001111100000110000110000000001100011000000000010001110000000001100001110000000110000011110000011000000001111111000; 
      9'd165: data <=256'b1111111111000000100000001100000000000000111000000000000011000000000000001100000000000111100000000001111111000000000011001111000000000000001111000000000000000110000000000000011100000000000000110000000000000011000011100001111100000111111111000000000111110000; 
      9'd166: data <=256'b0011111111111000111110000001110000000000000111000000000000111000000000001111000000000011111111100011111111111111011110000000001101100000000001100000000000011110000000000011100000000001111100000000001111000000001111110000000011110000000000001110000000000000; 
      9'd167: data <=256'b0000011111111110000111100000000001111100000000000111000000000000111000000000000011000000000000001100000000000000110000000000000011000000000000001110011111111110111011000000111111111100000001110111110000000011001111000000011100001111101111100000011111111100; 
      9'd168: data <=256'b0011111111111100011100000000110000000000000011100000000000001110000000000001110000000000111110000111111111110000011111111111100000010000000011100000000000000110000000000000011100000000000001110000000000001110110000001111111011111111111100001111111110000000; 
      9'd169: data <=256'b0000000000011111000000000111100000000001111000000000001100000000000011110000000000011000000000000011111100000000011111111000000011111000111000001110000001100000111000000110000011000000011000001100000011000000110000011000000011111111100000000011100000000000; 
      9'd170: data <=256'b0000000000000111000000000000111000000000000011100000000000011100000000000111110000000000111111000000000111011100000000111001110011111111000111001111100000011100000000000001100000000000000110000000000000111000000000000011100000000000001110000000000000111000; 
      9'd171: data <=256'b0000000000011111000000000111100000000001111000000000011111000000000011100000000000001110000000000011110000000000001110000110000001111011111111000111111111111110011111000000011001110000000011101111000000111100111111011111100000111111111000000000011100000000; 
      9'd172: data <=256'b0000000011111111000000011100000000000011100000000000001100000000000001110000000000000111000000000000011000000000000001100000000000000111000000000000011100000000000000111000000000000011100000000000001110000000011011111000000011111110000000001111100000000000; 
      9'd173: data <=256'b1111111111100000000000001110000000000000111000000000000011000000000000001100000000000001110000000000000111000000000000011000000000000001100000000000000110111111000000111111100011111111110000001111111110000000000000111000000000000001100000000000000110000000; 
      9'd174: data <=256'b0000111111111000011111000111110011111000001111101111000000000111111000000000000111000000000000111100000000000011100000000000001110000000000001101000000000001110100000000001100011000000000000001100000000000000111100000000000001111111100000000000010000000000; 
      9'd175: data <=256'b0000000000111110000000011110000000001111000000000000110000000000001110000000000001110000000000001100000000000000110000000000000011001111111110001111100000001100111000000000111101110000000000110011100000000011000111100000011100000111111111100000000001110000; 
      9'd176: data <=256'b0000000000011100000000001111100000000000111000000000001110000000000001110000000000001110000000000001110000000000001110000000000000110001111111100110011110000111011111100000001111110000000000111110000000001110111100000011110010111111111110000000011110000000; 
      9'd177: data <=256'b0000000000000000011111111111111111111111111111111100000000000000110000000000000011000000000000001101111110000000111111111111000000100000001111000000000000011110000000000000111000000000000111100110000000111100011111001111100000011111111000000000000000000000; 
      9'd178: data <=256'b0000000111000000000001111100000000001110011000000001100001100000011110000110000011100000011000001100000001100000100000000110000011110000011000000111111111111111000000000110000000000000011000000000000011100000000000001110000000000000111000000000000011000000; 
      9'd179: data <=256'b0001000001111111000110111111000000111111100000000111000000000000011000000000000011100000000000001100000000000000111111000000000011111111100000000000000111000000000000001100000000000000110000000000000011000000000000011100000000000111000000000000011000000000; 
      9'd180: data <=256'b0000001111111000000011110001100000111000000110000000000000011000000000000001100000000000001100000000000001110000000000000111000011000000111000001111111111111111000000001100000000000001110000000000000111000000000000011100000000000001110000000000000110000000; 
      9'd181: data <=256'b0000000001111111000000011110000000000011110000000000011100000000000011100000000000011110000000000001111110000000001111111110000001111000111100001111100001111000111100000011100011110000000110000011000000011000001110000011100000011111111100000000111000000000; 
      9'd182: data <=256'b0000111111000000000111111111100000111111001111100001100000000011000110000000011100001100000111000000111011111000000000111100000000000111110000000011111111000000011100000110000011100000011100001100000000110000110000001111000011111111110000000011111000000000; 
      9'd183: data <=256'b0000000111111110000011111100011000111000000001101110000000000110111110000000110000000000000110000000000001110000000000000110000000000001111111100000111100000111000111000000001100000000000000110000000000000011000000000000011100001111111111000000000001000000; 
      9'd184: data <=256'b0000011111111000000011110001111000011100000011100011100000111100001110001111100000111111111111110011111110000000011111000000000011111110000000001100011100000000110001111000000011100011100000000111000111000000000111001110000000001111111000000000001111100000; 
      9'd185: data <=256'b0000011111111110001111110000111011111000000111101000000001111000000000001110000000000111100000000001111000000000000111111111000000011111111111100000000000000111000000000000011100000000000011100000000000111100000001111111100011111111000000000011110000000000; 
      9'd186: data <=256'b0000000000011111000000000011111100000000001110110000000000111011000000000011101100000000001110110000000000111110000000000011111000000000001111000000000000111000000000000111100000000000111110000000001111011100000011110001110001111110000010001111000000000000; 
      9'd187: data <=256'b0001111111000000001110001110000001110000111000000110000001100000011000000110000001101100111000000111110011100000000000001100000000000001100000000000011110000000000011110000000011111110000000001111000000000000001111000000000000011111111111110000000011111000; 
      9'd188: data <=256'b0001111111110000001110000011110001110000000011101100000000000010110000000000001111000000000000111000000000000011110000000000001111000000000000111100000000000110011000000000110001110000000110001101110001110000110001111110000001110111100000000011111100000000; 
      9'd189: data <=256'b1111111111100000111111111111000000000000011110000000000001111000000000111111000000001111110000000001111110000000000011111100000000000011110000000000000111111000000000000011110000000000000111100000000000011110000001111111111100000111111111000000000011000000; 
      9'd190: data <=256'b0000111111110000000111000001111001110000001111111110000000111111111000000111111011100011111111101111111111111100001111111101110000000000000111000000000000011100000000000001110000000000001111000000000000111000111000001111000001111111111000000000111110000000; 
      9'd191: data <=256'b0000000000111000000000001111100000000000111100000000000011110000000000011110000000000011111000000000011111000000000111111100000011111101110000001100001110000000000000111000000000000011100000000000001110000000000000111101111001111111111111110001111111000000; 
      9'd192: data <=256'b1111111111111110000000000000011100000000000001110000000000001110000000000001111000000000001110000000000001110000000000001100000000000001110000000000011110000000000011111111100001111111111110000111100000000000111100000000000011000000000000001100000000000000; 
      9'd193: data <=256'b0000011111111100001111110000011101110000000000111110000000000111110000000001111011000000001111101111111111111110001111111100011000011111000001100000000000000111000000000000011100000000000001110100000000000111111100000000011001111111111111000000011111100000; 
      9'd194: data <=256'b0000111111110000001110000001100001110000000011001100000000001100110000000000110011110000001110001111100111110000011111111111111100011111110011100000000000001100000000000001110000000000001110000000000000110000000000000111000000000000111000000000000011000000; 
      9'd195: data <=256'b0001111111111110111111000001111111100000000000001110000000000011111100000001111101111000011111000011111111100000000011111000000000011111110000000011110111111000111100000011110011100000000011111111000000000111011110000000111100011111111111100000001111100000; 
      9'd196: data <=256'b0000111111111000001111000011110001110000000001101110000000000110110000000000001011000000000000111100000000000011111000000000001111100000000000111110000000000010111110000000001011100000000001101110000000011110011100000011100000111011111000000000111110000000; 
      9'd197: data <=256'b0000000000111000000000011111000011111111111100001111000001100000000000000110000000000000110000000000000011000000000000001100000000000001111111110011111111111100111111111100000001100001100000000000000111000000000000011100000000000000111000000000000001100000; 
      9'd198: data <=256'b0000011111111100001111111001111001111100000011101111100000000110111100000000011011110000000001111111000000000110111100000000111011100000000111101110000000011100111000000011110011100000011100001110000011110000011100011110000001111111110000000001111110000000; 
      9'd199: data <=256'b0011111111100000011100000111000011100000001100001111100000110000111111100111110011111111111111000111111111011100000000000000110000000000000011100000000000000110000000000000011100000000000001110000000000000111000000000000011111111111111111101000000111111100; 
      9'd200: data <=256'b0000000110000000000000111000000000000111000000000000011000000000000011000000000000011000000000000011100000000000001100000000000001110000000000001110000000011111110000000011011111000111111001111111111000001100011000000001110000000000001110000000000000110000; 
      9'd201: data <=256'b0000001111111110000111111110000001111100000000001110000000000000111100000000000001111100000000000000111111100000000000001111100000000000001111000000000000001111000000000000011100000000000000110000000000000111000110000111111000111111111110000001111110000000; 
      9'd202: data <=256'b0000000111111000000011111000000000011100000000000011100000000000011100000000000011100000000000001100000000000000110000000000000011000000000000001100000000111000110001111111111111111111000000110111110000000011011110000000111100011111111111000000111111000000; 
      9'd203: data <=256'b1111000000000000000111100000000000000110000000000000011100000000000001110000000000000111000000000000011000000000000001100000000000001100000000000001110000000000001110000000000000110000000000000111000000000011111000000000001111111111111111100011111100000000; 
      9'd204: data <=256'b0000000000111000000000001110000000000011100000000000111100000000000011000000000000111000000000000111000000000000111000000000000011000000000000101100000000001111110000000111111011100011111111000111111110111000000000000011100000000000001110000000000000011100; 
      9'd205: data <=256'b0000000001110000000000000111000000000000011100000000000001110000000000001111000000000000111000000000000111100000000000011110000000000011111000000000111111110000000111001111000011111000011100000000000001110000000000000011111100000001111111110000000011111100; 
      9'd206: data <=256'b0000011111100000000011001111000000000100001110000000000000111000000000000011100000000000011100000000000011100000000000011100000000000111100000000000111100000000001111000000000001111000000000001111000000000000110000000000000011111111111111110111111111111000; 
      9'd207: data <=256'b0000011111110000000011100111000000001000000110000001100000011000000110000001110000010000000110000000000000011000000000000011000000000000011100000000000011100000000000011100000000000111100000000000111100000000011111111111100011111111111111111100000000001100; 
      9'd208: data <=256'b0000011111111111000011110000000000000001110000000000000011000000000000001110000000000000011000000000000001110000000000000011000000000000001100000000000000111000000000000001100000000000000111000000000000011100111111110001110001111011111110000000000000100000; 
      9'd209: data <=256'b0000011000000011000111100001111100111111111111000110111111100000110000000000000011000000000000000111000000000000001110000000000000011100000000000000111000000000000001100000000000000110000000000000111000000000000111000000000011111000000000001111000000000000; 
      9'd210: data <=256'b0000001110000000000011111000000000011111000000000011110000000000011110000000000001110000000000001111000000000000111000000000000011100000000000001110000000000000111000000000011101110000001111100011111111111100000111111111110000000000011110000000000001110000; 
      9'd211: data <=256'b0000000000111111000000001111011100000000111011110000000111011100000000011111100000000001111100000000011111000000000011111110000001111111110000001110000011000000110000001100000011000000110000001100000111000000111100111000000001111111000000001111111000000000; 
      9'd212: data <=256'b0001111111111100111111100000111000000000000011100000000000111100000000000111000000000111111000000001110000000000000111000000000000011111111100000000000011111000000000000001111000000000000001110000000000001110000000000001110000000111111110001111111100000000; 
      9'd213: data <=256'b0000000001111110000000011110000000000011100000000000111100000000000111000000000000111000000000000111100000000000111100000000000011100000000000001111111111111100111110000001111011000000000001111110000000000011011100000000011100111111111111100000111111100000; 
      9'd214: data <=256'b0000110000000000000001000000000000001111000000000000011100000000000001111000000000000111100000000000011110000000000001111000000000000111110000000000001111000000000000111100000000000001110000000000000111100000000000011110000000000000111000000000000001110000; 
      9'd215: data <=256'b0000001111111000000001110011100000001110001110000000110000111000000011100011000000001111111100000000000011100000000000001100000000000001110000000000001110000000000001110000000000000110000000000000111000000000111111000000001111111111110001111100000111111111; 
      9'd216: data <=256'b0000001111110000000011110000000000001110000000000001100000000000001100000000000001110000000000000110000000000000111000000000000011100000000000001111111111111110111000000000011101110000000000110111000000001111001111000111110000011111111100000000001110000000; 
      9'd217: data <=256'b0000111111000000000111101110000001111100011000001110000001100000111111001110000000000000110000000000000011000000000000011000000000000011100000000000001100000000000001110000000000000110000000000000110000000000000111000000011100011111111111000000111100000000; 
      9'd218: data <=256'b0000000111111110000000110000011000000000000000110000100000000011000111100000001100111000000000110011000000000011011100000000001111100000000001101100000000000110110000000000110011000000000110001100000001110000110000001110000011110111100000000111111000000000; 
      9'd219: data <=256'b0000000000001111000000000001111000000000011110000000000011100000000000011100000000000011100000000000011100000000000011100000000011111100000000000011110000000000001111110000000001110011100000001110000111000000111000111100000011111111100000000011111000000000; 
      9'd220: data <=256'b0000000111111110000000111000011100000110000000110000110000000011000111000000001100111110000001110011100000000110001110000000111001111000000011000110000000111000111000000111100011000000111000001100000111000000110001111000000011111110000000000111110000000000; 
      9'd221: data <=256'b0000111111111000000000000011110000000000000011110000000000000011000000000000001100000000000000110000000000000111000000000000011000000000000111000000000000110000000000011110000000000011100000000000011000000000111111000000000011110000000110001111111111110000; 
      9'd222: data <=256'b1111111111111100111000000000111000000000000001110000000000000111000000000000111000000000001111000000000111110000000000111110000000000000111111000000000000001110000000000000111100000000000001110000000000000110011111000011111000111111111110000000111111100000; 
      9'd223: data <=256'b1111111100000000100000111100000000000001110000000000000011100000000000011100000000000001110000000000001110000000011111111111111100001111111111000001111000000000000111000000000000111100000000000011100000000000011100000000000001110000000000000111000000000000; 
      9'd224: data <=256'b0000111111111100000111000000111000111000000000110011100000000011000111000000001100001111000011100000001110111100011111111111100011100000001110001100000000001100111000000000111001110000000001100001100000000011000011110000011000000011111111100000000000011000; 
      9'd225: data <=256'b0111111111100000111100001110000000000000011100000000000000110000000000000111000000000000111000000000001111000000011111111000000011111111111000001111000011111100000000000000111000000000000001110000000000000111000000000001111100011100011111000000111111111000; 
      9'd226: data <=256'b0000110000000000000011000000000000011000000000000011100000000000001100000000000001110000000000000111000000000000111000000000011111100000000001101100000000011100111010111111110001111111101110000000000000111000000000000111000000000000011000000000000001100000; 
      9'd227: data <=256'b1111111000000000011111110000000000000011000000000000001100000000000000110000000000000011000000000000011000000000000001100111111101111111111111101111111000000000000001100000000000000110000000000000011000000000000001100000000000000111000000000000001100000000; 
      9'd228: data <=256'b0001111111100000111110000110000010000000011000000000000001100000000000001110000000111111110000000111111111111000001111000011110000000000000011100000000000000111000000000000001101100000000001111110000000011110110000000011110011111111111100000000010000000000; 
      9'd229: data <=256'b0000011111000000000001101110000000001100011000000000110000100000000011011011000000000101101000000000011100110000000000000110000000000000011000000000000001000000001111101100000001100111100000111100011110000111100011110000110011111111111111000000000011100000; 
      9'd230: data <=256'b0000000001111111000000001111011100000011100000110000011100000000000011100000000000011000000000000011100000000000011111110000000011111111111000001111000001110000110000000011000011000000011100001100000111100000110011111000000011111110000000000011000000000000; 
      9'd231: data <=256'b1111111111111000110000000011100000000000001110000000000001110000000000001111000000001111110000000001111000000000011110000000000001111000000000000001111111111000000000000011111100000000000001110000000000001111000000000111110000001111111000000001111100000000; 
      9'd232: data <=256'b0011111111111100011100000000000011100000000000001100000000000000111000000000000001111110000000000001111111100000000000000011100000000000000111100000000000000111000000000000001100000000000000110000000000000011000010000000011100001111111111100000001111111000; 
      9'd233: data <=256'b0000000111111110000000000000111100000000000011110000000000001111000000000001111000000000001111100000000000111000000000000111100000000001111110000000001111100000000001111100000000001111000000000011111000000000011111000000000011100000000000001000000000000000; 
      9'd234: data <=256'b0000000000000000000000000011111100000000111001110001111110000011001101100000001101100000000000110110000000000011010000000000001011000000000000101100000000000010100000000000011011000000000011001100000000011000011111110000000000001100000000000000000000000000; 
      9'd235: data <=256'b0000111111110000001111111111110001111000000011001111000000000110111000000000011011000000000001101100000000000111111000000000011111100000000001110110000000000011011100000000011101111000000001110011110000001110000111100011110000001111111110000000001111100000; 
      9'd236: data <=256'b0000000001111000000000000111100000000000011100000000000011110000000000001111000000000000111000000000000011100000000000011110000000000011110000000000001111000000000000111100000000000011100000000000111110000000000011110000000000011111100000000000111000000000; 
      9'd237: data <=256'b0000000011111110000000111100011100000110000001110000111000001110000111000011110000011100011100000000111111100000000001111000000000011111110000000111100011100000111000000110000011100000011000001100000011100000110000011100000011111111100000000001110000000000; 
      9'd238: data <=256'b0000000011110000000000111111000000000111000000000000111000000000000111000000000000111000000000000111000000100000111000001111110011000011111111101100011100000111110001100000001111001100000001111110011000001111111001100001110001111111111110000001111111100000; 
      9'd239: data <=256'b0000000011111100000000111101110000000111000011000000011000001100000001100011110000000111111011000000001111011100000000000001100000000000001110110000000001110011001111000110001101111111110000111100001111111111100011111111111011111100000000001111000000000000; 
      9'd240: data <=256'b0001111111110000001110000011000000110000000110000010000000110000000000000111000000000000111000000000001111000000000001110000000000001100000000000011100000000000011100000000000011100000000000001100000000000111110000111111111111111111111000000111110000000000; 
      9'd241: data <=256'b1111111100000000110001111110000000000001111110000000000000111000000000000001110000000000000111000000000000011100000000000011100000000000011110000000000011110000000001111110000000000111100000000001111000000000111111000001111111111111000111001111111111100000; 
      9'd242: data <=256'b0011111000000000001100110000000000110001100000000001100010000000000111111000000000000111100000001110011111100000001111100110000000000000001100000000000000111000000000000000110000000000000011100000000000000011000000000000001100001111010111100000011111111100; 
      9'd243: data <=256'b0111111111111100111000000000110001000000000111000000000000111000000000000111100000000000111000000000001111000000000001110000000000011110000000000011100000000000011100000000000011100000000000001100000000000000100000000000000011111111111111110011111111000000; 
      9'd244: data <=256'b0011111111000000111100001110000010000000011000000000000001100000000000000110000000000001111000000100011110000000111111111110000000000000011111000000000000001110000000000000011000000000000000110000000000000011011100000000001111111111111111110000111111111100; 
      9'd245: data <=256'b0001111111111110011110000000001111100000000111111110000000111100011100001111000000111111111000000000111111000000000111001111000001111000001111101110000000001110110000000000011011000000000001111100000000000110011110000011111000011111111100000000001110000000; 
      9'd246: data <=256'b0001111111111110011110000000111111100000000000111110000000000111111000000000011101111111100111100111111111111100000111111111000000000000011100000000000011100000000000001110000000000001110000000000001111000000000000111000000000000111000000000000011000000000; 
      9'd247: data <=256'b0001100000000000001110000000000001110000000000001110000000000000111000000000000011000000000000001100000000000000110000000000011111100000000011111110000001111110011110011111110000111111110111000000000000011100000000000001110000000000000011100000000000000111; 
      9'd248: data <=256'b0000000001111100000000000000011000000000000000110000011100000011000111110000001100111000000000110111000000000011011000000000001011000000000000101100000000000110100000000000110010000000000110001000000000110000110000001110000001111111100000000011111000000000; 
      9'd249: data <=256'b1111111111110000110000001111100010000000001110000000000000111000000000000111000000000011111000000000011110000000000011100000000000111100000000000011100000000000111100000000000011100000000000001100000000000000111000011111111111111111111000000011111110000000; 
      9'd250: data <=256'b0000000000111110000000000111100000000000111100000000001111100000000001111100000000001111000000000001111000000000000111000001000000111111111111000111111111111111011110000000011111110000000011111111000000011110111110001111110000111111111100000011111111000000; 
      9'd251: data <=256'b0000000001111110000000000100001100000000000000110000000000000011000000000000011000000000000011100000000000011000000000000011000000000001111000000000001110000000000111100000000001110000000000001100000000000000110000000000000011110000000000000011111111111100; 
      9'd252: data <=256'b0111111111000000111100001110000000000000001100000000000000011000010000000000100011000000000011001100000000001110110000000000011011000000000001111100000000000011011000000000001101100000000000110011000000000110000111000000111000001111111110000000001111110000; 
      9'd253: data <=256'b0000110000000000000011000000000000011100000000000011100000000000001110000000000000110000000000000111000000001111011000000001111111100000000111111100000000111110110000000011110011111111111110000000000000111000000000000011100000000000000111000000000000000110; 
      9'd254: data <=256'b0001111111111111000110010000000100000000000000000001100000000000001100000000000001100000000000001110000000000000111111100000000011111111100000000000000111000000000000001100000000000000110000000000001110000000000001110000000001111110000000000011100000000000; 
      9'd255: data <=256'b1111111111100000100011111111100000000000000111000000000000111000000000000111100000000011111000000001111110000000001111000000000001111111000000000011111111111100000000000001111100000000000000110000000000000111000000001111111011111111111110000011110000000000; 
      9'd256: data <=256'b0001111111110000001110000011100000110000000110000010000000011100000000000001100000110000000110000001111111111100000000000000010000000000000001100000000000000011000000000000001100000000000000110000000000001110100000000011110011100000111100001111111111000000; 
      9'd257: data <=256'b0000000000011111000000000111001100000000111000000000000111000000000001111000000000000110000000000001110000000000000110000000000001111001100000000110001111000000111011101100000011111000110000001111000111000000111000111000000011111111000000000011110000000000; 
      9'd258: data <=256'b0000110000000000000111000000000001111000000000001111000000000000111000000000000011000000000000001100000000000000111100000000000001111111111111110000000000000111000000000001111000000000001110000000000000111000000000000011000000000000001100000000000000010000; 
      9'd259: data <=256'b0000001111110000000000111110000000000011110000000000001111000000000000111000000000000111100000000000110111000000000111011100000001111000110000001110000011010000110000111111111111111111110000111111000011000000000000001110000000000000111000000000000011100000; 
      9'd260: data <=256'b0000011111100000000001101110000011001100011000001110110001100000001111111100000000011000000000000011100000000000001100000000000000110000000000000011000000000000011111111111111111110000000000001011100000000000001100000000000000011000000000000001100000000000; 
      9'd261: data <=256'b0000000011111110000111111000111011111100000111000000000001110000000000001111000000000001110000000000000110000000000000110000000000000111000000000011111111111111000111000000000000011000000000000001100000000000001110000000000000110000000000000001000000000000; 
      9'd262: data <=256'b0011111111110000011100000011110000000000000011100000000000001110000000000001110000000000011110000000111111100000011111110000000001111111111100000000000000111110000000000000011000000000000000110000000000000111000000000000111011111111111111001111111110000000; 
      9'd263: data <=256'b0000011111111111000111100000001101110000000000011110000000000011110000000000111011000000001111101111111111111100000000000000110000000000000011000000000000001100000000000000110000000000000011000001000000001100000111000000110000001111111111000000000011111000; 
      9'd264: data <=256'b0111000000000000001100000000000001110000000000000110000000000000011000000000000011100000000000001100000000000000110000000000110011000000000111001100000000011100110000000011110011100000111111000111111111101100000011100000111000000000000011100000000000000111; 
      9'd265: data <=256'b0000001111111110000000111111011000000111100000110000011100000011000001100000011100000110000011100000111001111100000011101110000000001111110000000001111110000000011111100000000011001110000000001000110000000000110011000000000011011100000000000111100000000000; 
      9'd266: data <=256'b0000011111111100000011110000111000011100000001100011100000000011001100000000001101110000000000110111000000000011111000000000001111100000000001111111000000000110111100000000111011110000000011001111100000011100011111000111100001111111111100000011111111000000; 
      9'd267: data <=256'b0000000011111110000000000000011100001100000000110000110000000110000011000011110000001100111000000000111111000000001111100000000011110111000000001100001100000000110000011000000011000001110000000110000011100000001110000110000000001111111000000000000110000000; 
      9'd268: data <=256'b1110000000000111011100000001111000111111111111000110011111110000011000000111000001100000111000001100000111000000100000111000000011000111111000001111111111000000000011000000000000011100000000000011100000000000011100000000000001110000000000000110000000000000; 
      9'd269: data <=256'b0000011111111100001111100001111001111000000011100110000000011100111110000011110011111111111100001000001111100000100011111111000000011110011110000001110000011100000110000001111000011000000011100001100000000111000011100000111000001111111111000000001111110000; 
      9'd270: data <=256'b0000000000011100000000000001110000000000001111000000000001111100000000000111100000000000111111000000000011110000000000011111000000000011111000000000001111000000000001111100000000001111100000000001111100000000001111110000000000111100000000000001000000000000; 
      9'd271: data <=256'b0000000000111111000000111111000000111111000000000011000000000000011100000000000011100000000000001100000011000000110111111111000011111100000111100000000000000111000000000000011100000000000001110000000000001110000000000111110011100111111000000111111100000000; 
      9'd272: data <=256'b0000000111111111000011111000000000111100000000000011000000000000000110000000000000001100000000000000111000000000000001110000000000000001100000000000000011100000000000001111000000000000001100000000000000111000100000000011100011110001111100000111111111100000; 
      9'd273: data <=256'b0011100000000000001111000000000000001111000001110000111111111111000011000011100000001100111000000000110111000000000000111000000000000111000000001111111111110000111111111111000000011100000000000011100000000000001100000000000000110000000000000011100000000000; 
      9'd274: data <=256'b0000000000000111000000000001111100000000011110000000000011100000000000111100000000000011000000000000111100000000000111000000000000111001111100000111111111111000011110000001110011100000000111001100000000111000100000000111000011111111110000000000110000000000; 
      9'd275: data <=256'b0000000000010000000000000011000000000001101100000000001110111000000001110011000000001100001100000011100000110111011000000011110011100000111110001111111111100000111100000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000; 
      9'd276: data <=256'b0000111111111110001111000000011101100000000000110110000000000011011000000000001100110000000011100011000000111100001111011110000000001111100000000011111110000000111100001110000011000000011100001100000000111000111000000011000000110000011100000001111111000000; 
      9'd277: data <=256'b0000000011000000000000011100000000000011100000000000011110000000000011100000000000011100000001110111100000001111011100000000111111100000000011111111111000011111001111111111111000000011111111000000000000111000000000000011100000000000011110000000000000110000; 
      9'd278: data <=256'b0000000111111110000000110000011111100000000000110011000000000111000111100000111000000111001110000000000111110000000000011110000000000111001100000000110000011000001110000001110001110000000111000110000000011000111000000110000011111111110000000011111000000000; 
      9'd279: data <=256'b0000000011100000000000001110000000000001111000000000000111000000000001111110000000001110111000000001110011100000001100001110000011100000011000000000000001100000000000000110000000000000001100000000000000110000000000000011000000001111111111100000000111111111; 
      9'd280: data <=256'b0000000000000111000000000000111100000000001111000000000001111000000000011110000000000111111000000000111111000000001111111000000011111111000000000000111000000000000111000000000000111000000000000111000000000000011100000000000001100000000000000111000000000000; 
      9'd281: data <=256'b0000000000000011000000000000001100000000000000110000000000000111000000000000111100000000000011110000000000111111000000000011011000000000011001100000000111000110000000111000011000000111000001100001110000000110001100000000011111100000000001111000000000000000; 
      9'd282: data <=256'b0000001111110000000011110000000000011100000000000011110000000000011110000000000011110000000000001110000000000000111000000000000011111111111110001111111111111100111100000000111011111000000011111111110000001111000011100000111100001111111111110000000011111000; 
      9'd283: data <=256'b0011111111111110001110000011111100000000000001110000000000111110000000011111100000000011110000000000001111100000000000001111000000000000001110000000000000011100000000000000110000000000000011100000000000001110111100000001111011111111111111000000011111100000; 
      9'd284: data <=256'b0000000011111111001111111111000000110000000000000000000000000000110000000000000011111110000000001111111110000000111000111100000010000000111000000000000001100000000000000110000000000000001000000000000001100000001000000110000000111111111000000001111110000000; 
      9'd285: data <=256'b0000000001111111000000000000111000000000001111000000000011100000000000001111000000000000001110000000000000011100000000000000110000000000000011000000000000011100000000000011000000000000011100000000011111100000000111110000000011111000000000001110000000000000; 
      9'd286: data <=256'b1000000000000000110000000011000001100000001100000011111111110000000011111100000000000001100000000000000110000000000000011000000000000011000000000000111111111111000000110000001100000011000000000000001110000000000000011000000000000001100000000000000011000000; 
      9'd287: data <=256'b0000000000000111000000000000111100000000000111000000000000111100000000000111100000000011111100000000111101110000111111000111000011110000011000000000000011100000000000011100000000000011100000000000011100000000000001110000000000000110000000000000011000000000; 
      9'd288: data <=256'b0011000000000000001100000000000001100000000000000110000000000000011000000011000011100000001100001100000000110000110000000011000011000000001100001100000011111111111111111111000000000000001100000000000000110000000000000010000000000000001000000000000000100000; 
      9'd289: data <=256'b0000000000011111000000000111100000000000111000000000001111000000000001110000000000000110000000000001110000000000001110000000000001110000000000001111111111111110111110000000111011110000000001101110000000111110111110001111100000111111111000000000010000000000; 
      9'd290: data <=256'b0000000000000011000000000000011100011110111111100000011111011000000000000001100000000000001100000000000001110000000000000110000011111111111111001111111111111111000000011100000000000001100000000000001110000000000000111000000000000011000000000000001100000000; 
      9'd291: data <=256'b1111111111111000111111100001110000000000001110000000000111110000000001111100000000111110000000000111100000000000000111111100000000000000111111100000000000001111000000000000111100000000000111100000000001111000000001111110000000111111000000001111000000000000; 
      9'd292: data <=256'b0000001111111111000000110000000000000110000000000000111000000000000111000000000000111111111110000011111111111110001110000000111000000000000011100000000000011110000000000011110000000000001110001111100111111000111101111110000011111111100000000011111000000000; 
      9'd293: data <=256'b1111111111100000000000001111100000000000011110000000000011110000000000111100000000011110000000000001111111110000000000000111000000000000000111000000000000000110000000000000011000000000000000110000000000000111000000000001111010001111111111001111111000000000; 
      9'd294: data <=256'b0000000111111111000011111000011100001100000001110000000000001110000000000001110000000000001110000000000011100000000000111100000000000111100000000000111000000000001111000000000001110000000000001110000000000000111000000000000011111111111100000111111000000000; 
      9'd295: data <=256'b0001110000000000001110000000000001110000000000001111000000000100111000000000111011100000000011111100000000011111111000011111111111111111111111100000000000011110000000000001111000000000000111100000000000011110000000000001110000000000000111000000000000011100; 
      9'd296: data <=256'b0111111111000000110000001100000010000000110000000000000011000000000000001100000000000001110000000000001110000000000000111000000000000011000000000000111100000000000011100000000000011100000000000011100000000111111110001111111001111111111000000000111100000000; 
      9'd297: data <=256'b0000000011000000000000001100000011111111110000000000000011000000000000011100000000000001110000000000000111000000000000011000000000001111111111110111111110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000; 
      9'd298: data <=256'b0000000000001111000001111111111000001111000000000011110000000000000110000000000000011000000000000001110000000000000011000000000000001100000000001100110000000000110011000000000011001110000000001100110000000000110011000000000001111000000000000011000000000000; 
      9'd299: data <=256'b0001111111111000000110000001110000100000000111000110000001111000011000011110000001111111100000000111111100000000111101111000000011000001111000001000000001111000110000000001111001100000000001110111000000000011000111000000001100001111001111110000001111111100; 
      9'd300: data <=256'b0000100000000000000110000000000000011000000000000011000000000000011000000000000001000000000000001100000000000000110000000000000011000000000001001100000000001100111000000111110001111111110011000000111100001100000000000000110000000000000011100000000000000111; 
      9'd301: data <=256'b0011100000000011011110000000111101111000000111100111000011111000111111111110000010000001110000000000001110000000000001110000000011100111111110001111111111000000010110000000000001111000000000000111000000000000111000000000000011000000000000001000000000000000; 
      9'd302: data <=256'b0000011111111111000111111000000000001110000000000000110000000000000011000000000000011100000000000001100000000000000111110000000000111111110000000001000011100000000000000111000000000000001100000000000000110000000000000111000011111111111000000111110000000000; 
      9'd303: data <=256'b1111111110000000110000011100000000000000111000000000000001110000000000000011000000000000001100000000000000110000000000000011000000000000011000000000000011100000000000011000000000000011100000000000001100000000000000111000000000000001111111110000000011111110; 
      9'd304: data <=256'b0000000000011000000000000011000000000000011100000000000011100000000000111100000000000111000000000001110000000111001110000000110111110000000011111100000000001111111110000000111100111111101111100000000111111100000000000000110000000000000011100000000000001110; 
      9'd305: data <=256'b0011111111111110011111111000011111111100011111111111000001111110111000001111110011111111111100001111111111111000000000000011100000000000001111000000000000011100000000000011110000000000001110000000000001111000000000001111000000000011110000000000111100000000; 
      9'd306: data <=256'b1111111000000000011011111000000000000001110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000001100000000000111110000000000111111111111100000011000000000000011100000000000001100000000000001110000000000000110000000000; 
      9'd307: data <=256'b0000110000000000000111000000000000011000000000000011100000000110011000000000011001100000000011001100000000011000110000000001100011000000001100001111100011111111011111111110000000000000110000000000000110000000000000010000000000000011000000000000011000000000; 
      9'd308: data <=256'b0000000001111100000000111110111000001110000001110011110000001111011000000001111111011000001111111101111111110111111111111000011100000000000001110000000000000011000000000000001100000000000000110000000000000011000000000000111101111111111111110001000000000000; 
      9'd309: data <=256'b0000011111100000000011100011100001111100001011001101100000000110110110000000011011011000000000111000100000000011100010000000001110001100000000111000000000000011110000000000011111000000000001100110000000001100011110000011110000011111111000000000111111000000; 
      9'd310: data <=256'b1111111111110000110000000111100010000000001110000000000001111000000000001111000000000011111000000000011100000000000011100000000000111100000000000111000000000000111000000000000011000000000000001100000000000000111111111111111101111111110000000000010000000000; 
      9'd311: data <=256'b0000000111111111000001111110000011000000000000001100000000000000110000000000000011000000000000001111110000000000000011100000000000000111000000000000001110000000000000011000000000000011100000000000001110000000011001110000000001111110000000000001110000000000; 
      9'd312: data <=256'b0000000111111000000001111000111000000110000001110000011000000111000001100000111100000111111111100000011111111111000001111100001100000000000000110000000000000011000000000000001100000000000000111110000000000011011111000000001100011111111111110000000011111100; 
      9'd313: data <=256'b1111111100000000110000111000000010000011100000001100001110000000000000111000000000000111000000000000111111111000000000000001110000000000000011100000000000000111000000000000011100000000000001110000000000001110000000000001110000000011111100000000001111100000; 
      9'd314: data <=256'b0000000000001111000000000000111100000000000111100000000000111110000000000111110000000000111110000000011111111000000111110011110011111100001111000000000000111100000000000011110000000000011111000000000000111000000000000011111100000000001111110000000000000100; 
      9'd315: data <=256'b0000001111111100000001111000111000011110000001110011110000000111011110000000001111111000000000111111000000000011111100000000001111000000000000111100000000000111111000000000111011100000000011100110000000011100011110001111100000111111111000000001111110000000; 
      9'd316: data <=256'b0000000111111100000001111100111100001110000000110001110000000000001110000000000000110000000000000111000000000000111000000000000011100000000000001110000011111100111000111101111111100111000001111110011000000111111000110000111101111011001111000011111111111000; 
      9'd317: data <=256'b0000001111111111000001110000011100001110000001110001110000001110000111000001110000001100001110000000110111110000000011111111000001111111000000001110001110000000110000111000000011000001110000001110000011100000011100000110000000111111111000000000011110000000; 
      9'd318: data <=256'b0000000000111110100000000110011011110000011111100111111111111000000000000110000000000000011000000000000001100000000000011111111100000001111111110000000111100000000000001111000000000000011100000000000000110000000000000011000000000000001110000000000000011000; 
      9'd319: data <=256'b0000000000001111000000000000111000000000000011100000000000001110000000000000111000000000000111100000000000011110000000000111111000000001111011101000011110001110111111110000111001000000000011100000000000001110000000000000111000000000000011100000000000001100; 
      9'd320: data <=256'b0000000001110000000000000111000000000000011100000000000011110000000000001110000000000001110000000000001111000000000001111000000000000111100000000000111100000000000011100000000000011110000000000001110000000000000111000000000000011100000000000000111100000000; 
      9'd321: data <=256'b0000000000000111000000000000111100000000000011100000000000111100000000011111110000000011100011000001111100001100011110000000110011100000000011000000000000001100000000000000110000000000000011000000000000001100000000000000111000000000000011100000000000000100; 
      9'd322: data <=256'b1111111111110000000000000111000000000001111000000000111110000000000111100000000000111100000000000001111100000000000001111111100000000000011111100000000000000111000000000000011100000000000011100000000000111000000000011111000000011111100000000001100000000000; 
      9'd323: data <=256'b0000111111111110000111000000111100111000000001110011100000000011001100000000011100111000000001110001110000001111000011100000110000000111111111000000111111111000111111001111000011000000001110001100000000011100111000000000110001111111111111000000111111111000; 
      9'd324: data <=256'b0001100000000000000110000000000000110000000000000111000000000000011100000000000111110000000000111100000000000011110000000000011111000000000011101100000000001110110000000011111011100000111011100111111111000110000000000000011100000000000001110000000000000011; 
      9'd325: data <=256'b0001111111111100001111100001111000111100000011100111000000001110011100000000011111100000000001111110000000000111110000000000011111000000000001111110000000000111111000000000011111110000000011110111100000011110001111111111110000011111111100000000001111000000; 
      9'd326: data <=256'b0000000000011000000000000001100000000000001110000000000001111000000000001111000000000011101100000000011101110000000011000110000000111000011000000110000001111111110000011111100011111111110000001111110011100000000000001110000000000000111000000000000001000000; 
      9'd327: data <=256'b0000011110000000000011100000000000011100000000000001100000000000001100000000000001110000000000000110000000000000111000000000011111000000000001101100000000001110110000000000111011100000111011000111111110001110000000000000111000000000000001100000000000000010; 
      9'd328: data <=256'b0000000011111000000000111100000000001111100000000000110000000000011111000000000001110000000000001110001111111100111011111111111011111100000001111111100000000111111000000000011111100000000011101110000000011100111110000111100000111111111000000000111111000000; 
      9'd329: data <=256'b0000000000011100000000000001110000000000000110000000000000111000000000000111100000000000110110000000001110011000000001100001100000011100000110000011000000011000111000000001100000000000000110000000000000011000000000000001101100000000011111110000000001110000; 
      9'd330: data <=256'b0000000111111111000000111000000000000111000000000000000000000000001111000000000001110000000000001111111100000000000000111100000000000001111000000000000011110000000000000011100000000000001110000000000000111000000100001111100000011111111000000000011110000000; 
      9'd331: data <=256'b0000000111111111000001111000011100001110000000000011110000000000001110000000000001111000000000001110000000000000111000000000000011000001111100001100011111111000110111111111110011111000000111001111000000111100111000000011100011111111111110000011111111000000; 
      9'd332: data <=256'b0011111111111110111000000000001011000000000000111110000000001111111000000001100000110011111100000111111111100000011011100000000011100011100000001110000111100000011100000110000000110000001110000011100000011100000011100000111000000111100011100000000111111100; 
      9'd333: data <=256'b0000000000001111000000000000111100000000000111100000000000011100000000000011110000000000011111000000000011101100000000011000110000000111100011000000111000001100000111000000111000111000000011101111111111111110111111111111111000000000000011100000000000000110; 
      9'd334: data <=256'b0000111111100000000111111100000000111000000000000111000000000000111000000000000011011111111000001111110111111100000000000000111000000000000001110000000000000011000000000000001100000000000001110000000000001110001000000000110000111000111110000001111111000000; 
      9'd335: data <=256'b0011111111111110111110000000011101110000000000110111100000000011011111000000011100111110011111100000111111111110000000111110111100000000000001110000000000000111000000000000011100000000000001111111000000001111111111000011111000011111111110000000001111000000; 
      9'd336: data <=256'b0111111111000000111000001110000001000000111000000000000011100000000000001110000000000001110000000000001110000000000001110000000000001110000000000001110000000000001110000000000001110000000000001110000000000000110000000000000011111111111111110111111111000000; 
      9'd337: data <=256'b0000111111100000000111000011000000011100001100000001110000110000000011100011000000000111011000000000001111111000000011111100000001111111111000001110000001110000110000000001110011000000000011000110000000000111001110000000001100001111000001110000001111111110; 
      9'd338: data <=256'b0000000000000011000000000000011100000000000001100000000000011110000000000001111000000000001111000000000011101100000000011100110000000011100011000000111100001100000111000000110000111000000011000111000000001100110000000000110011000000000001000000000000000100; 
      9'd339: data <=256'b0000001111100000000011110000000000011110000000000011100000000000011100000000000011100000000000001110000000000011011111111111111100011111000111100000000000111000000000001110000000000001110000000000001110000000000001110000000000000111000000000000001111100000; 
      9'd340: data <=256'b0000000000110000000000000110000000000000110000000000000110000000000000110000000000001110000000000001100000000000001110000000000001110000000000001110000001111111110011111100011011111100000011001111000000001100000000000011100000000000011100000000000011100000; 
      9'd341: data <=256'b0111111111100000111000000111100010000000000111000000000000001100000000000000110000000000000111000000000000111000000000111111000000000111111000000000000111111100000000000001111100000000000000110000000000000011000000000000011100000011111111100000000101100000; 
      9'd342: data <=256'b0000011100011110001111000000001111000000000000011100000000000011011100000000011100111000000111000000111101111000011111111111000011111111111110001111000000110000100000000001100010000000000110001000000000011000000000000011000000111111111000000000110000000000; 
      9'd343: data <=256'b0000111111100000000110000111000000000000011100000000000011110000000000011100000000000111100000000000111111110000000000000011100000000000000111100000000000000110000000000000011100000000000001110000000000011110000000000111110011111111111100000001100000000000; 
      9'd344: data <=256'b0000000111111110000000010000011000000000000000110000000000000011000000000000011100000000000111000000011111111000000001111101110000000000000011100000000000000111000000000000001100000000000000110000000000000111000000000000111011001001111111001111111111000000; 
      9'd345: data <=256'b0000001111111100000001111001110000011111000011100011111000000111001111000000011101111000000000111111100000000011111100000000001111100000000000111110000000000011111000000000001111100000000001111111000000001110101100000001110010011110001110001000111111110000; 
      9'd346: data <=256'b0000011111000000000000011100000000000011111000000000000111100000000000011110000000000001111000000000000111100000000000011110000000000001111000000000000111100000000000111110000000000011111000000000001111000000000000111100000000000011110000000000001110000000; 
      9'd347: data <=256'b0000000111111000000000111111110000001111000111000001110000011000001110000011100001110000011100001110000011100000110000011100000011000001100000001100001100000000000001100000000000001110000000000000111000000000000001111100111100000001111111100000000001111000; 
      9'd348: data <=256'b0000000000000011000000000000011100000000001111100000000001111100000000111111100000011111011100000111100011100000111000011100000011000011100000001110011111111000011111111111000000001100000000000001110000000000001110000000000001110000000000000111000000000000; 
      9'd349: data <=256'b0000001111111100000001111000110000001110000001100001110000000110001110000000001101110000000000111100000000000011110000000000001111000000000000111110000000000011011000000000011101110000000011100011100000001100001111000001110000001111111110000000011111100000; 
      9'd350: data <=256'b0000011110000000000001111000000000001111110000000000110111000000000111011100000000111000110000000111100011000000011000001100000011100000111000001100000011100000110000001111111111111111111110000111111111100000000000000110000000000000011000000000000001100000; 
      9'd351: data <=256'b0001111111111100001110000000111001110000000000100110000000001110011100000111110000111111111100000111111111100000111001110000000011000001111000001100000000111000011000000000110001110000000011110001110000000011000001110000001100000011111111110000000001111100; 
      9'd352: data <=256'b0000000011111110000011111111000000111100000000000111000000000000111000000000000011100000000000001111111111000000000000111111000000000000011111000000000000001110000000000000011100111110000000110111100000000111011100000000111101111111111111100000111111110000; 
      9'd353: data <=256'b0000111111111111001111110000000001110000000000001110000000000000110000000000000011011100000000001111111110000000111000111110000011100000111100000000000000111000000000000001100000000000000110001111000000111000111100000111000001111111111000000000011110000000; 
      9'd354: data <=256'b0000000001111111000000001110001100000001110000010000000110000001000000011000001100000001100001100000000110011100000000011111000011111111111000001100000010000000100000001100000010000000110000001100000001000000011000000110000000111111110000000000001100000000; 
      9'd355: data <=256'b0000000000000111000000000001111000000000000111000000000001111100000000001111110000000011110110000000011100011000000111100011100001110000011100001110000001110000100000001110000000000000111000000000000011100000000000001100000000000001111000000000000011100000; 
      9'd356: data <=256'b0111111111111000111000000001110011100000000011100110000000000011011100000000001100111000000011110001111111111100000001111000000000011111111111100011111110000000111100011000000011000001100000001100000011000000110000011100000011111111110000000001111100000000; 
      9'd357: data <=256'b0011111100000000011111111000000001100001111000000010000001100000000011111111000000000111100100000000000000010000000000000001000000000000001100000000000001100000000000011110000000000011000000000111111000000000111000000000000011111111111111000000000000000111; 
      9'd358: data <=256'b0000111111100000111111111110000011111100000000000111000000000000011100000000000001111111000000000111111111100000011111111111000011110000001111000110000000001110000000000000011100000000000000110000000000000011000110000000111100011111111111000000111111111000; 
      9'd359: data <=256'b0000000111111110000000111000001100000011000000110000011000000011000001100000011000000111000111000000011111111000000000011111100000000111100111000001111000011100001100000000111001100000000011101100000000111100100000001111100011110111111000000111111100000000; 
      9'd360: data <=256'b0000000000011111000000001111000000000011111000000011111110000000001110000000000001100000000000001110000000000000110000000000000011100000000000000111111111100000000000000011000000000000001100000000000011100000001100111100000011111111000000000111100000000000; 
      9'd361: data <=256'b0011111111000000111110011110000011000000011100000000000011110000000000011110000000000111100000000011111000000000111111100000000000111111111000000000000011111000000000000001111000000000000001110000000000000111000000000000111100111111111111100000011111100000; 
      9'd362: data <=256'b0000001111111100000011111100111100001110000000110000110000000011011101110000001111000001111111111111000011111100011111111111000000000000001100000000000000110000000000000011100000000000001110000000000000111000000000000001100000000000000110000000000000011000; 
      9'd363: data <=256'b0000110000000000000011000000000000001100000000000001100000000000001110000000000000110000000000000110000000000000011000000000010011100000000001101100000000000110110000000000011011000111111111101111111111101111000000000000011100000000000001100000000000000110; 
      9'd364: data <=256'b0000000111111110000001111000100000001111000000000001111000000000001111000000000001111000000000000111000000000000111100000000000011110000000000001110011111110000110111111111110011111100000111101111100000001111011110000000111000111111111111100001111111111000; 
      9'd365: data <=256'b1111111111110000000000000011100000000000001110000000000001111000000000001111000000000000111000000000001111000000000000111100000000001111000000000001110000000000001111000000000000111000000000000111000000000000111000000001111101111111111110000111111110000000; 
      9'd366: data <=256'b0000000011100000000000001100000000000001110000000000001111000000000001111100000000001100110000000011110011000000011100001100000011100000110000000000000110000000000000011000000000000001100000000000000110000000000001110000000001111111100011110001111111111110; 
      9'd367: data <=256'b0000000011111000000000000000100000000000000110000000000000011000000000000011100000000000011100000000000011100000000000011000000000000111100000000000111000000000000111000000000000111000000000001111000000000000110000000001111111111111111110000001100000000000; 
      9'd368: data <=256'b0000000000111111000000000111001100000000110000110000000110000011000001110000001100001110000001100000110000000110000110000000110011111000000111001110000000011000111000000011100011000000011100001100000011100000111000111000000011111111100000000011111000000000; 
      9'd369: data <=256'b0011111111111111001110001111111101111000000000000111000000000000011100000000000001110000000000000111000000000000001100000000000000011111100000000000001111000000000000001111000000000000011100000000000001110000000010001111000011111111111000001111111110000000; 
      9'd370: data <=256'b0000001111000000000001110110000000000110011000000000011101100000000000110110000000000000011000000000000001100000000000001110000000000000110000000000000111000001000000111000001100001111000000111111111000000110111111110000111011100011111111000000000011111000; 
      9'd371: data <=256'b0001111111000000011110001110000011000000011110001100000000111000000000000011100000000000001110000000000000111000000000001111000000000011111000000000111100000000011111100000000011100000000000001110000000000111111000000011111111111111111110100000001000000000; 
      9'd372: data <=256'b0000000011110000000000001111000000000001111100000000000011110000000000011110000000000001111000000000001111000000000001111100000000001111100000000000111100000000000011110000000000011110000000000001111000000000000111000000000000011100000000000001100000000000; 
      9'd373: data <=256'b0000000000001110000000000001110000000000001110000000000011100000000000011100000000000011100000000000111000000000000011000000000000111100000000110011100000000111011000000000111111100000011111111100111111100111111111100000011000000000000001100000000000000010; 
      9'd374: data <=256'b1111111111111111000000000000011100000000000011100000000000011110000000000011100000000000001100000000000011110000000011001100000000001111111111000000011111100000000001110000000000001110000000000001111000000000000111100000000000011110000000000000110000000000; 
      9'd375: data <=256'b0001111111111111011111000000000011000000000000001100000000000000110000000000000011000000000000001101111100000000111110110000000011110001100000000000000110000000000000011000000000000001100000000000000100000000000010110000000000001011000000000000111000000000; 
      9'd376: data <=256'b0000111111100000000000000011100000000000000110000000000000011000000000000111100000000000111000000001111111000000000111111100000000000000011111000000000000000110000000000000001100000000000000110000000000001110000000000011110001011111111100001111111100000000; 
      9'd377: data <=256'b0000111111111100111111000000111010000000000011100000000000001110000000000001110000000001111110000011111111111000001111110001110000011100000011110000000000000011000000000000001100000000000001110000000000001111111100000001111001111111111110000000000110000000; 
      9'd378: data <=256'b0000000000011111000000001111111000000001111000000000001110000000000011110000000000111100000000000011100000000000011100000000000011100000000000001100011111100000111111111110000011111000011100001110000001100000111000001110000001111111110000000001111100000000; 
      9'd379: data <=256'b0000000000111100000000001111110000000111110111000000111000011000000111000001100001110000000110001110000000011100110000000001100011100000000110000111000000011000001111111111111100000000011110000000000000011000000000000001110000000000000011000000000000001100; 
      9'd380: data <=256'b0111111111000000000111111111000000111000001110000111000000011100011000000000011011000000000001111100000000000011110000000000001111000000000000111100000000000011111000000000001101111000000001110001111000001110000011111111110000000000111100000000000000000000; 
      9'd381: data <=256'b0000000011110000000000011111000000000001111100000000001111110000000011110111000000001110110000000001110011000000000110001100000001110000110000001111000111001111110001111111111111111111111111001100000110000000000000111000000000000011100000000000000110000000; 
      9'd382: data <=256'b0011111111111000001100000001111000000000000011100000000000000110000000000000111100000000000011100000000000011100000000000111100000000011111000000000111100000000001111000000000001111000000000001110000000011111111100011111100001111111111000000000111000000000; 
      9'd383: data <=256'b0111111111111100001000000001111100000000000000110000000000000111000000000000111000000000001111000000000001110000000000011110000000000111100000000000110000000000011110000000000001100000000000001100000000000000110000000000000011111100000000000000110000000000; 
      9'd384: data <=256'b1100000000111110110000000111111111100000011111100111111111111100000000011110000000000001110000000000000111000000000000011000000000011111110000000000111111111100000000111000000000000011000000000000001100000000000000110000000000000011100000000000000100000000; 
      9'd385: data <=256'b0001111111110000001100000001110000110000000011100011000000000110000110000000011000111110000111100001111111111000000000111100000000001111111110000111111000111000111000000000111011000000000001111100000000000011111000000000001101111000000001110000111111111110; 
      9'd386: data <=256'b0111111111111111011000000000000011000000000000001100000000000000111111110000000001111111111000000000000001110000000000000011000000000000000110000000000000011000000000000001100000000000000110000000000001110000000000001110000000000111100000000001111100000000; 
      9'd387: data <=256'b0000111111000000111111111100000011111100000000000110000000000000111000000000000011000000000000001100000000000000111111111110000011111111111111000000000000001110000000000000011000000000000001110000000000000111000000111000111000000011111111000000000011111000; 
      9'd388: data <=256'b0000011111110000000011110011100000111100001110000010000000110000000000000111000000000000111000000000000111000000000000110000000000001110000000000000110000000000001110000000000001110000000000001110000000111111110000011111111111111111111001101111100000000000; 
      9'd389: data <=256'b0000011111111100011111100001111100111110000001110011111000000111000111000000111000011110000111000000111000111000000011111111000000000111110000000000011111000000000111111100000000011011110000000111001110000000111001111000000011111110000000001111000000000000; 
      9'd390: data <=256'b0111100000000000111111111111000011111111111111111110000000000000111000000000000011000000000000001110000000000000111100000000000001111111111000000000000011110000000000000011100000000000000110000000000000111000000111111111000001111111110000000111100000000000; 
      9'd391: data <=256'b0000000000001111000000000001111100000000001111100000000001111110000000011110110000000011100011000000111100011000000011000001100001111000001111001111111111111000111111111111100000000000001100000000000000110000000000000011000000000000001110000000000000011000; 
      9'd392: data <=256'b0000011111111111001101000000000000100100000000000011100000000000000110000000000000001100000000000000111000000000000001100000000000000011000000000000001100000000100000011000000010000001100000001100000011000000011100001100000000011111100000000000011110000000; 
      9'd393: data <=256'b0000000000111100000000001111000000000001110000000000011110000000000011100000000000011110000000000011100111111000001111111000111001111100000000110111000000000011111100000000001111110000000000111111000000001110111110000001110011011111111110001000001111000000; 
      9'd394: data <=256'b1111111000000000110011110000000011000011000000000000001100000000000000111000000000000011000000000000001100000000000011111111111111111111110000001100001100000000000000110000000000000011000000000000001100000000000000100000000000000110000000000000010000000000; 
      9'd395: data <=256'b0111111110000000000000011000000000000000110000000000000010000000000000011000000000000011100000000000011100000000000011100000000000111100000000000111000000000000111000000000000011000000000000001100000000000000111110000000011001111111111111110000110011111111; 
      9'd396: data <=256'b0000000111111110000011110000001100111000000000010111000000000011111000000000001111100000000111101111000001111100011111111111100000011111111110000000000000111000000000000011100000000000001100000000000000110000111000000011000011111111111100000000001111100000; 
      9'd397: data <=256'b0001111111111111111111111111000011100000000000001110000000000000110000000000000011000000000000001100000000000000111000000000000001111000000000000001110000000000000011110000000000000011100000000000000111000000011000001100000001111111110000000000111110000000; 
      9'd398: data <=256'b0000000000011100000000000111110000000000111110000000000011110000000000011111000000000011111000000000001111000000000001111000000000000111100000000000111100000000000111110000000000011110000000000001111000000000001111000000000000011110000000000000001000000000; 
      9'd399: data <=256'b0000001111111111000111111110011100011000000001110001110000001110000011000001100000001110011110000000011111100000000001111100000000000011100000000000011110000000000111111000000000011001100000000111101110000000111001110000000011111110000000001111100000000000; 
      9'd400: data <=256'b0000011111110000000111110011100000011100000000000001110000000000000011111111111100000111111100110000000000000111000000000000011000000000000011100000000000001110000000000000110000000000000011000000000000011100000000000001110011111111111111001000111111111000; 
      9'd401: data <=256'b0011111111100000011110011111000011100000111100001110000001111000111000000011100011100000001111000111000001111100001111111111111000000111000011100000000000000110000000000000011100000000000001110000000000000111000000000000111100000111111111100000011111100000; 
      9'd402: data <=256'b0001100000000000000110000000000000111000110000000011000011000000011100001100000011100000100000001100000110001111110000011111111111111111111111101111000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000; 
      9'd403: data <=256'b0000001111111100000001111110110000001111110001100001111100001111000111101111111000011101111101100011111111000110001111110000110001111110000011000111100000001100011100000011100011100000001100001111000011110000111100011100000010111111100000000001111000000000; 
      9'd404: data <=256'b0000000000011111000000000111000000000001111000000000001111000000000001111000000000001110000000000011110000000000001110000000000001111000000000001111011111111100111111100000111011111100000001101110111000001110111000000001110001111111111110000000011100000000; 
      9'd405: data <=256'b0000011111111110001111100000011000000000000001110000000000001110000000000001110000000000001100000000000111100000000001110000000000011100000000000111100000000000110000000000000010000000000000001100000000000000111000000000000001111111001111110001111111111000; 
      9'd406: data <=256'b0000000000000011000000000000011100000000000001100000000000001110000000000000110000000000000111000000000000111000000000000111000000000000011100000000000011110000000000111110000000000110011000000000111001100000000111000110000011111000011000001110000000000000; 
      9'd407: data <=256'b0000000011111110000000111000010000001110000000000001100000000000001110000000000001110000000000001110000000000000111000000000000011100011111111101100111110111111110011100000111011101110000000101111100000000110011110000000110000111110011110000000111111100000; 
      9'd408: data <=256'b0000000011111000000000001001100000000000000110000000000000110000000000000111000000000000111000000000000111000000000000111000000000000111000000000000111000000000111111000000001111110000000001111111100000001110001110000011110000011111111110000000111111100000; 
      9'd409: data <=256'b0001111111111110001111000000011001110000000001111110000000111111110000000111111011111000111111100111111111111110000000110000111000000000000011100000000000000111000000000000011100000000000001100000000000011110000011100011110000001111111110000000001111100000; 
      9'd410: data <=256'b0000011111111100000001100001111000001110000001100001110000000011000110000000001100110000000000110111000000000011011000000000001111000000000000101100000000000110110000000000110011000000000011001110000000111000011110001111000000111111111000000000001100000000; 
      9'd411: data <=256'b0000000111111000000001111001110000000110000110000000111001111000000011101110000000000111110000000000111111000000001111001111000001110000001111000000000000001110000000000000011101100000000000111100000000000111111000000000011001111111111111100001111111110000; 
      9'd412: data <=256'b0000111111111111000110000000001100111000000000000111000000000000011000000000000001100000000000001111111111110000000000000011100000000000000110000000000000011000000000000000100000000000000110000000000000111000000000001111000010000011110000001111111110000000; 
      9'd413: data <=256'b0001111111111110111111111001111111111000000111111111000000011111111110000011111011000000001111001111111111111000000111110110000000000000111000000000000111000000000000111000000000000111000000000000011100000000000011100000000000001110000000000000111000000000; 
      9'd414: data <=256'b0000000011111110000000011110111100000011100000110000011100000011000001110000001100000111000011110000001110011100000000111111110000000111111100000001110011100000011100001111000011100000001110001100000000011000111000000001110001110000001110000001111111110000; 
      9'd415: data <=256'b0000001111111100000001110000011000001110000001100000110000000011001110000000001101110000000000110111000000000011111000000000001111100000000000111100000000000110110000000000011011000000000001101110000000011100011100000011100001111111111100000001111111100000; 
      9'd416: data <=256'b0000111111111000001111000001100000100000000110000000000001111000000000000110000000000000110000000000011111000000000011100000000000011110000000000111110000000000011100000000000011100000000000001110000000000000111000000000000011111110000000000011111111111111; 
      9'd417: data <=256'b0000001111100000000011111111100000111110001111100111100000001110011100000000011111100000000000111110000000000011110000000000001111000000000000111100000000000111111000000000011111100000000011100111100000011100001111100111100000001111111100000000001110000000; 
      9'd418: data <=256'b1111111111000000110000111111000000000000001100000000000001110000000000011110000000111111100000000011111111110000000000001111100000000000001111100000000000000111000000000000011000000000000011100000000000011110000000000111100001111111111000000011111000000000; 
      9'd419: data <=256'b0000000111000000000000011100000011100011110000000111101111000000000111110000000000000011000000000000001000000000000000101111111111111111111111111110001000000000100000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000; 
      9'd420: data <=256'b0000000000111000000000000111000000000000111000000000000111000000000000111000000000000111000000000000111000000000000111000001100000111000001100000111000000111000111000000011100011000000001110001100011111111111111111111001110011111000000011000000000000000100; 
      9'd421: data <=256'b0000000111111110000000111111110000001111110000000001110000000000001111000000000000111000000000000011111111111000001111100011110000010000000011100000000000000110000000000000011100000000000001111110000000000111111000000000111111111111111111100000011111110000; 
      9'd422: data <=256'b0011111111100000111100000111100011000000000111001000000000001110110000000000011000000000000001100000011000001110000001111100110000000111111110000000000000011100000000000000011000000000000000110001100000000011000111000000001100001111110111110000000111111100; 
      9'd423: data <=256'b0000000000000111000000000001110000000000001100000000000011100000000000111000000000000110000000000000110000000000000110000000000000111000000000000110000111111100011001110000011011011100000001001100000000011100110000000011100011110011111000000011111110000000; 
      9'd424: data <=256'b0000011111111000000111111011111000111100000001110111000000000011011110000000111100111100111111100000111111110000111111111100000011100011110000001110000011100000111000001111000001110000001110000011100000011100000111100001110000000111111111000000000011110000; 
      9'd425: data <=256'b0000000000011111000000000111110000000001111100000000001111000000000001110000000000001110000000000001110000000000001110001111100001110111111111100111111000000110111110000000011011111000000001101111000000001110111111000011110011101111111100000111111111000000; 
      9'd426: data <=256'b0001111111111100011110000011111100000000000001110000000000000111000000000001111000000011111110000011111110000000000111111100000000000001111110000000000000011110000000000000011100000000000000110000000000000011000000000000111111000000111111001111111111000000; 
      9'd427: data <=256'b0000000111111110000011111100011100111100000000110111000000000111011100000000111001111111111111000011111111111000000001100111100000000000111100000000000111000000000000111100000000001111000000000001111000000000011111000000000011110000000000001100000000000000; 
      9'd428: data <=256'b0000000000111111000000001111001100000011111001110000011100001110000001100001110000001100011110000000110011100000000111111100000000011111110000000011100011100000011100001100000011100000110000001100000111000000100001111000000011001110000000000111110000000000; 
      9'd429: data <=256'b0000001110000000000000111111000000011111111110000111100011110000111100000111100011000000011111001100000011111100111000011100111001111111100001110000000000000011000000000000001100000000000000110000000000001111011100000001111001111111111111000000011111100000; 
      9'd430: data <=256'b1111111111111111011000000000000001000000000000000100000000000000110000000000000011000000000000000110000000000000011000111110000001111111111110000000000000001100000000000000110000000000000111000000000000011000110000000011100011111111111100000111111110000000; 
      9'd431: data <=256'b1111111111111110111111111110000010000000000000001100000000000000011111111111110001110000000001100100000000000011000000000000000100000000000000110000000000000110000000000000010000000000000011000000000000111000000000000010000000000000111000000000000110000000; 
      9'd432: data <=256'b0000000001111110000000001110001100000000110000110000000000000011000000000000011100000000000011100000000000011110000000000011100000000011111110000000111110000000111111100000000011111100000000000000111100000000000000111000000000000011111100000000000011110000; 
      9'd433: data <=256'b0000001111111110000011110000001100011110000000110011110000001111001111111111111000111000100000000111000000000000011000000000000011100000000000001110000000000000111000000000000011100000000000001110000000000000111000000000000011111000000000001111100000000000; 
      9'd434: data <=256'b0000011111111110000111100000001100111000000000110111000000000110011000000001111001110000011100000111111111100000111111111111110011111000000000001101110000000000110011100000000011100111000000000110011100000000011100111000000000111111100000000001111110000000; 
      9'd435: data <=256'b0000000111100000000000111110000000000111100000000000111000000000001111100000011001111000000011100111000000001110111100000000111011111100000111100111111111111111000111111111111100000000111100000000000011100000000000011110000000000011100000000000011100000000; 
      9'd436: data <=256'b0000000000000111000000000000011000000000000011100000000000001100000000000000110000000000001111000000000000111100000000000111100000000001111110000000001100111000001111100011100001111000001110001100000000111000000000000011100000000000001111000000000000111000; 
      9'd437: data <=256'b0001111111110000001111001111111000111000000011110011110000000111000011100000111100000111111111110000011111110000000111111100000001111100111100001111000001111000111000000001110011100000000011101111110000001110111111111111111001111111111111100000011111111000; 
      9'd438: data <=256'b0000000001111111000111111110001111111000000001101100000000000110000000000000110000000000000011000000000000011000000000000001000000000001111100000000001111111100000000001110000000000000110000000000000011000000000000011100000000000001100000000000000110000000; 
      9'd439: data <=256'b0000011111111111000000000000111000000000000111000000000000111000000000001111000000000000110000000000011110000000111111111110000011111111111110000001110000000000001110000000000001111000000000000111000000000000111000000000000011000000000000001000000000000000; 
      9'd440: data <=256'b0011111111111110000110000000110000011000000000000011100000000000001100000000000000111111111100000111000001111100001100000000111000000000000001100000000000000111000000000000001111100000000000111100000000000111111100000000111000111111111111000000111111110000; 
      9'd441: data <=256'b0111111111111111011111111111100001100000000000000110000000000000011000000000000001100111111110000111111000011100001110000000111000000000000001100000000000000110000000000000011000000000000001110000000000000111000000000000011111111111111111100000011111111100; 
      9'd442: data <=256'b0111111111110000111110000011000001110000000000000110000000000000011000000000000001111000000000000011111111000000000000111111110000000000000011100000000000000111000000000000011100000000000001110010000000000111011111000000111000111100001111000000111111110000; 
      9'd443: data <=256'b1111111111100000111000001111000011000011111000000000011100000000000001100000000000000111000000000000001111000000000000001110000000000000011110000000000000011100000000000000111000000000000001110000000000000011000000000000011100001111111111100000000111100000; 
      9'd444: data <=256'b0000000000000000000011111111100000011100000011100011100000000111011000000000111111100000000000011100000000000011110000000000011111000000000001101100000000001100110000000011100011100000011100001110000011100000011111111000000000111111000000000000000000000000; 
      9'd445: data <=256'b0011111000000000001101110000000000110011000000000011100110000000001110011000000000011111100000000000111110000001000000011000001101111001100001111111111110000110110001111000111011000011110011001100001111101100111111110111110001111110000111000001100000001100; 
      9'd446: data <=256'b0001111111110000011111000111110011100000000111101101111000011110101110000000111100111000000001110011000000001111001110000001111100011110011111110000111111110011000000000000001100000000000000110000000000000111000000000000111000000111111111000000000111110000; 
      9'd447: data <=256'b0000001111111100000011110000111000011100000001110001100000000011001100000001111101110000000111100111000000111110011100000011100000111111111111000001111110001100000000000000111000000000000011110000000000000111000000000000011111111111111111101110000000000000; 
      9'd448: data <=256'b1110000000000000011110000000000000001100000000000000010000000000000001100000000000000100000000000000110000000000000011000001111100011111111110010001100000000000001100000000000000110000000000000110000000000000011000000000000001100000000000000110000000000000; 
      9'd449: data <=256'b0000000001111000000000011111000000000001111000000000001111100000000000111110000000000011110000000000011111000000000001110000000000001111000000000000111000000000000011100000000000011110000000000011110000000000001110000000000000011000000000000000111000000000; 
      9'd450: data <=256'b0000001111000000000000111100000000000111110000000000011011000000000011101100000000011100111000000011100001100000001100000111000001110000011100000110000000110000111000000011100011100000001110001110000000111111011100011111100001111111110111000000000000001100; 
      9'd451: data <=256'b0011111111100000111111001110000010000000011100000000000001110000000000000110000000000000011000000000000001100000000000000110000000000000011000000000001111100000000000011111111100000000111000000000000011100000000000001110000000000000110000000000000011000000; 
      9'd452: data <=256'b0000000011111111000000111000000100000011000000010000001000000011000000100000000000000011000000000000000111111000001111111111000011111101100000001000000010000000100000001000000011000000100000000110000010000000001000001000000000001111100000000000011100000000; 
      9'd453: data <=256'b0111110000000000111111100000000011000111100000001100001110000000111000011000000011111001100000000011110011000000000000001100000000000001110000000000000111000000000000111000000000001111000000000111111000000000001111111000000000000111111111110000000000011100; 
      9'd454: data <=256'b0111111100000000000000111000000000000001100000000000011110000000000111100000000001111000000000001111100000000000001111111000000000000001111110000000000000011110000000000000011000000000000001110000000000001111000000000001110011111111111110000011111110000000; 
      9'd455: data <=256'b0000111111111100000111111001111001111100000001110111000000000011111000000000001111100000000000111100000000000011110000000000001111000000000000111100000000000110110000000000111011100000000111001110000000111000011100001111000000111111110000000001111110000000; 
      9'd456: data <=256'b0000000000000111000000000000011100000000000001110000000000000111000000000000111000000000000011100000000000011110000000000001110000000000001111000000000001111100000000011111110000000001100111000000011110011100000011100000000001111100000000001110000000000000; 
      9'd457: data <=256'b0000011111111111000000000011100000000000011100000000000011000000000000011000000000000011100000000000001100000000000000100000000011110110000000001111110000001111011111111111111000011000000000000001100000000000000110000000000000110000000000000011000000000000; 
      9'd458: data <=256'b0000000111100000000000011110000000000011111000000000001111100000000000111100000000000111110000000000011110000000000011111000000000001111000000000000111100000000000011110000000000001110000000000000111000000000000011100000000000000111000000000000000110000000; 
      9'd459: data <=256'b0000000000111111000000000111100000000001111000000000001111000000000001111000000000001110000000000011110000000000001110000000000001111000000000001111001111111000111111110011100011111100001110001111100011110000111000111100000011111111100000000111110000000000; 
      9'd460: data <=256'b0111111110000000111000111100000010000001111000000000000111000000000000111100000000000111100000000000111100000000000011100000000000011100000000000001110000000000000111000000000000001110000000000000111100000000000001111000000000000011111111110000000011111110; 
      9'd461: data <=256'b0000000111110000000000111011000000000011001100000000001100110000000000110011000000000011011000000000000001100000000000001100000000000001110000000000001110000000000000110000000000001110000000010011111110000011011100111110011011110000111111101100000000000000; 
      9'd462: data <=256'b0000000000000111000000000000011100000000000001110000000000000111000000000000011000000000000011100000000000001110000000000011111000000000001111100000000011100110000000001100011000000011110001100000011100000110001111100000000011111000000000001100000000000000; 
      9'd463: data <=256'b0111111110000000110000001100000010000000110000000000000011000000000000011100000000000011100000000000111000000000000011111000000000000001111000000000000000111000000000000000111000000000000001110000000000000011000011000000011100001100011111100000011111110000; 
      9'd464: data <=256'b0000000000000000000000011111100000000111110111000000111100001110000111110000011000111111000001110011110000000011011110000000001101110000000000111111100000000111111010000000111011100000001111001111111111110000001111111100000000000000000000000000000000000000; 
      9'd465: data <=256'b0000000001111100000001111110000100011111000000110001100000000111000110000001111000111000011110000001101111100000000111111000000000011110000000000011111000000000011111100000000011100111000000001100001110000000111000011000000000111101100000000000111110000000; 
      9'd466: data <=256'b0000000011111100000001111100111000011110000011110011100000000111111100000000111111000000001111101100000011111100111111111101110001111110000111000000000000011100000000000011100000000000001110000000000001110000000000001111000000000111111000000000001100000000; 
      9'd467: data <=256'b0000001111111100000001111000111000000000000011100000000000011110000000000001111000000000011111000000000011111000000000111110000000001111100000000011111000000000011111000000000011110000000000001110000000000000111000000000000011111111111111110000010010000000; 
      9'd468: data <=256'b0011111111100000000111111111110000000000000111100000000000001110000000000001111000000000001110000001111111110000000111111111000000000001111111100000000000001111000000000000011100000000000011110000000000111110111100011111100011111111110000000000100000000000; 
      9'd469: data <=256'b0000111111111000000111000100110000111000000011100011000000000110011000000000001011100000000000111110000000000011110000000000001111000000000000111100000000000011110000000000001111100000000000111110000000001110011110000011111000111111111110000000111000000000; 
      9'd470: data <=256'b1111111111100000110000000000000011000000000011111000000000011110110000011111100011000011110000001111111100000000011111000000000001111000000000001111110000000000110011100000000011000111100000001100000111000000011100011100000000011111110000000000011110000000; 
      9'd471: data <=256'b0000000000000000000111100000000000111111111100000111110000111100111000000000111011100000000001101110000000000111110000000000001111000000000000111110000000000011011000000000011101110000000011100011110000111100000111111111100000000111111000000000000000000000; 
      9'd472: data <=256'b0000000000000111000000000000011100000000000011110000000000011110000000000011111000000000011111100000000011111100000000011101110000000111110111000001111100011100001111000011110011111000001110000000000000111000000000000011100000000000001110000000000000110000; 
      9'd473: data <=256'b0111111111100000111100000111000000000000011100000000000001100000000000011110000000000011100000000000111000000000000111111111000000011100011111100000000000000111000000000000001100000000000001110000000000001111000000000011110000000001111100000000001111000000; 
      9'd474: data <=256'b0011111111111111000000000000011100000000000011100000000000011110000000000011110000000000011100000000111111111000111111111111000011000111100000000000111100000000000111100000000000111100000000000011100000000000011100000000000011110000000000001110000000000000; 
      9'd475: data <=256'b0111111111111100111100000000110000000000000011000000000000011000000000000011100000000000111100000000011111111000000011110001111000000000000011100000000000000111000000000000011100000000000001110000000000001110000000000011110001110011111110000111111110000000; 
      9'd476: data <=256'b0000001111111100000011111000111000111100000001110111111000000011111011100000011111000110000011101000011100011100000000110011100000000011111100000000001111100000000000111000000000001111100000000001111110000000001110111000000000111111000000000000110000000000; 
      9'd477: data <=256'b0000000000111111000000000111000000000011111000000000111100000000000011100000000000111100000000000011100000000000011100000000000011110001111111001110001100011100111001100001110011100000000110001110000000111000111000001111000001111111110000000011111100000000; 
      9'd478: data <=256'b0000000000111000000000000011100000000000001100000000000001110000000000001111000000000001111100000000001111110000000011100110000000011100011000001111100001100000110000000110000000000000011000000000000001100000000001101110111100000111111111110000000111000000; 
      9'd479: data <=256'b0000000000011111000000000111100000000000011110000000000011110000000000111110000000000011110000000000011111000000000011111000000000011111000000000011111011111000011110111111110001111111100111101111001111111110111100001111110011111111111110000111111110000000; 
      9'd480: data <=256'b0000000000000111000000000000111000000000000111000000000001111100000000000111110000000001110111000000001110011100000001110001100000111110000110001111000000011000100000000011100000000000001110000000000000011000000000000001100000000000000111000000000000001100; 
      9'd481: data <=256'b0001111111100000000111000111000000010000001100000000000000110000000000000111000000000000110000000000001110000000000000110000000000011110000000000011100000000000011100000000000011100000000000001100000000000000110000000000000011111111111111110001111100000000; 
      9'd482: data <=256'b0000000000011100000110000111110001111111111100000111000011100000111000001100000011100000110000000000000111000000000000011000000000000011100011110011111111111110000001111000000000000011000000000000001100000000000000110000000000000011100000000000001110000000; 
      9'd483: data <=256'b0000000000111110000000001111100000000001111000000000011110000000000011110000000000011110000000000011100000000000011100000000000011111111111111101111111000001111111110000000011111110000000011111111100000011110111111001111100011111111111000000111111110000000; 
      9'd484: data <=256'b0000000000000111000000000000111100000000000111100000000000111100000000000111100000000000111100000000001111100000000000111100000000011111100000001111111110000000111100110000000000000111000000000000011010000000000011111000000000001111000000000000011000000000; 
      9'd485: data <=256'b1111111110000000111110111000000000000001100000000000000110000000000000011000000000000011000000000000001100011111000001101111100001111111111000000111111000000000000011000000000000011000000000000001100000000000001100000000000000111000000000000001100000000000; 
      9'd486: data <=256'b1111111110000000011111111111100000000000001111000000000000011100000000000011110000000001111110000000111111100000011111110000000011111111111000000000000111111000000000000011111000000000000011110000000000001110000000000000111000000000111111000000000011110000; 
      9'd487: data <=256'b0011111111111000011000000001110001100000000001110110000000000011011100000000011100110000000001100001110000111100000011001111000000001111100000000111111100000000111000011000000011000001100000001000000011000000110000001100000001110000110000000011111110000000; 
      9'd488: data <=256'b0011000000000000011000000000000001100000000000000110000000000000111000000000000011000000000000001100000000001100110000000000011011000000000011101100000000001110111100001111111001111111100011100001100000001110000000000000011000000000000001110000000000000011; 
      9'd489: data <=256'b0000000011110000111111111111000011111111110000000000001110000000000000111000000000000011100000000000001100000000000001110000000000111111111111110111111111000000011111100000000000111110000000000001111000000000000011100000000000001110000000000000111000000000; 
      9'd490: data <=256'b0000111111100000000111111111000000111000000111000110000000001100110000000000011011000000000000101000000000000011100000000000001111000000000000110110000000000011011000000000011100110000000001100011100000001100000111100111100000001111111100000000000000000000; 
      9'd491: data <=256'b0001111111110000001110000011100001110000000111100100000000000110110000000000011011000000000000111010000000000011111000000000001111100000000000110110000000000011011000000000011001100000000001000110000000001100001110000111100000011111111000000000111110000000; 
      9'd492: data <=256'b1111111111100000111111111000000011110000000000001100000000000000011110000000000000011110000000000000011100000000000000011100000000000000111100000000000000011100000000000000111000000000000001100000110000000011000001110000000100000011101000110000000001111110; 
      9'd493: data <=256'b0011111110000000011100111100000011100000110000000100000011000000011000011100000000000011100000000000001110000000000000111111100000000000000111100000000000000110000000000000001111111000000000111110000000000110111110000001111000111111111110000000001110000000; 
      default: data<=256'd0;
    endcase 
  end 
endmodule 
