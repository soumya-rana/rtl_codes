`timescale 1ns/1ps
///////////////////////////////////////////////////////////////////////////////
// Company: Indian Institute of Science, Bengaluru
// Engineer: Soumya Kanta Rana
//
// Create Date: 14.11.2021
// Module Name: hidden layer calculator
// Project Name: ELM engine
// Target Devices: xc7a200tfbg484-2
//
////////////////////////////////////////////////////////////////////////////////
module input_to_hidden (input [255:0] img,
  input clk,
  input set,
  output reg signed [31:0] hidden_node,
  output reg [12:0] node_index,
  output reg multiplier_en);
  
  wire signed [15:0] weight;                             // takes the weight values generated by LFSR
  reg [8:0] counter;                                     // iteration variable that keeps count of input node
  reg [255:0] input_layer;                               // stores the image provided as input (input nodes)
  reg signed [31:0] ans;                                 // register where hidden node value is calculated
  lfsr RAND(clk, set, weight);                           // instantiate LFSR for generating weights

  parameter HIDDEN_NODES=13'd3000;
  assign img_bit=input_layer[8'd255-counter];            // value of current input node

  always @ (posedge clk) begin
    if (set) begin                                       // if set is high
      input_layer<=img;                                  // read input image and store in input_layer
      counter<=9'd0;                                     // reset iteration counter to 0
      ans<=32'd0;                                        // reset ans to 0
      hidden_node<=32'd0;                                // reset output to 0
      node_index<=13'd0;                                 // reset node_index to 0 (the node whose value is being calculated)
      multiplier_en<=1'b0;
    end
    else if ((counter != 9'd256)&(img_bit)) begin        // if all 256 input nodes are not covered and the input node value is 1
      ans<=ans+weight;                                   // add weight value to ans
      counter<=counter+1'b1;                             // increment iteration counter
      multiplier_en<=(counter==9'd1)?1'b1:1'b0;          // disable the multiplier of next stage from reading data
    end
    else if ((counter != 9'd256)&(~img_bit)) begin       // if all 256 input nodes are not covered and the input node value is 0
      counter<=counter+1'b1;                             // increment iteration counter (no addition)
      multiplier_en<=1'b0;
    end
    else if ((counter == 9'd256)&(node_index!=HIDDEN_NODES)) begin                    // if all 256 input nodes are covered
      hidden_node<=ans[31]?32'd0:ans;                    // assign RelU(ans) to output hidden_node
      node_index<=node_index+1'b1;                       // increment node index (the value denotes which hidden_node value is present at output)
      counter<=9'd1;                                     // reset iteration counter to 1
      ans[14:0]<=(input_layer[8'd255])?weight[14:0]:15'd0;     // set answer to weight times 1st input layer
      ans[31:15]<=(input_layer[8'd255])?{17{weight[15]}}:17'd0;// perform sign extension (if ans needs to be set to weight value
      multiplier_en<=1'b1;                                // enable the multiplier of next stage
    end
  end

endmodule
