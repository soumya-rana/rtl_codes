///////////////////////////////////////////////////////////////////////////////
// Company: Indian Institute of Science, Bengaluru 
// Engineer: Soumya Kanta Rana 
//
// Create Date: 17.11.2021
// Module Name: images ROM answers
// Project Name: ELM engine
// Target Devices: xc7a200tfbg484-2
//
////////////////////////////////////////////////////////////////////////////////
module test_images_answers(input [8:0] addr,  output reg [9:0] data);
  always @ (addr) begin 
     case(addr)
      9'd1: data <=10'b0000001000; 
      9'd2: data <=10'b0001000000; 
      9'd3: data <=10'b0000000010; 
      9'd4: data <=10'b0000001000; 
      9'd5: data <=10'b0100000000; 
      9'd6: data <=10'b0100000000; 
      9'd7: data <=10'b0010000000; 
      9'd8: data <=10'b0000100000; 
      9'd9: data <=10'b0000000001; 
      9'd10: data <=10'b0000100000; 
      9'd11: data <=10'b0100000000; 
      9'd12: data <=10'b0010000000; 
      9'd13: data <=10'b1000000000; 
      9'd14: data <=10'b0001000000; 
      9'd15: data <=10'b0000001000; 
      9'd16: data <=10'b0000000010; 
      9'd17: data <=10'b0000100000; 
      9'd18: data <=10'b0000000010; 
      9'd19: data <=10'b0000000100; 
      9'd20: data <=10'b0000001000; 
      9'd21: data <=10'b0100000000; 
      9'd22: data <=10'b0000000001; 
      9'd23: data <=10'b0000000010; 
      9'd24: data <=10'b0000000001; 
      9'd25: data <=10'b0001000000; 
      9'd26: data <=10'b0000010000; 
      9'd27: data <=10'b1000000000; 
      9'd28: data <=10'b0010000000; 
      9'd29: data <=10'b0000010000; 
      9'd30: data <=10'b0000000100; 
      9'd31: data <=10'b0000010000; 
      9'd32: data <=10'b0000000100; 
      9'd33: data <=10'b0001000000; 
      9'd34: data <=10'b1000000000; 
      9'd35: data <=10'b0000000010; 
      9'd36: data <=10'b1000000000; 
      9'd37: data <=10'b0000000001; 
      9'd38: data <=10'b0000010000; 
      9'd39: data <=10'b0000000001; 
      9'd40: data <=10'b0000010000; 
      9'd41: data <=10'b0100000000; 
      9'd42: data <=10'b0000000100; 
      9'd43: data <=10'b0000010000; 
      9'd44: data <=10'b1000000000; 
      9'd45: data <=10'b0001000000; 
      9'd46: data <=10'b0000100000; 
      9'd47: data <=10'b0001000000; 
      9'd48: data <=10'b0001000000; 
      9'd49: data <=10'b0000100000; 
      9'd50: data <=10'b0001000000; 
      9'd51: data <=10'b0010000000; 
      9'd52: data <=10'b0000000100; 
      9'd53: data <=10'b0000001000; 
      9'd54: data <=10'b0000000001; 
      9'd55: data <=10'b0100000000; 
      9'd56: data <=10'b0001000000; 
      9'd57: data <=10'b1000000000; 
      9'd58: data <=10'b1000000000; 
      9'd59: data <=10'b0000001000; 
      9'd60: data <=10'b0000010000; 
      9'd61: data <=10'b0000000100; 
      9'd62: data <=10'b0000001000; 
      9'd63: data <=10'b0000010000; 
      9'd64: data <=10'b0100000000; 
      9'd65: data <=10'b0000000100; 
      9'd66: data <=10'b0000000001; 
      9'd67: data <=10'b0000010000; 
      9'd68: data <=10'b0010000000; 
      9'd69: data <=10'b0000001000; 
      9'd70: data <=10'b0000000100; 
      9'd71: data <=10'b0000000010; 
      9'd72: data <=10'b0000000001; 
      9'd73: data <=10'b0100000000; 
      9'd74: data <=10'b0000010000; 
      9'd75: data <=10'b0001000000; 
      9'd76: data <=10'b0000000010; 
      9'd77: data <=10'b0001000000; 
      9'd78: data <=10'b0000001000; 
      9'd79: data <=10'b0000010000; 
      9'd80: data <=10'b1000000000; 
      9'd81: data <=10'b0000100000; 
      9'd82: data <=10'b0001000000; 
      9'd83: data <=10'b1000000000; 
      9'd84: data <=10'b0001000000; 
      9'd85: data <=10'b0000100000; 
      9'd86: data <=10'b1000000000; 
      9'd87: data <=10'b0000000001; 
      9'd88: data <=10'b0100000000; 
      9'd89: data <=10'b0000100000; 
      9'd90: data <=10'b0001000000; 
      9'd91: data <=10'b0000100000; 
      9'd92: data <=10'b0000010000; 
      9'd93: data <=10'b0000100000; 
      9'd94: data <=10'b0001000000; 
      9'd95: data <=10'b0000000100; 
      9'd96: data <=10'b0000000001; 
      9'd97: data <=10'b1000000000; 
      9'd98: data <=10'b0000000100; 
      9'd99: data <=10'b0000000100; 
      9'd100: data <=10'b0000000100; 
      9'd101: data <=10'b0000100000; 
      9'd102: data <=10'b0000001000; 
      9'd103: data <=10'b0000000001; 
      9'd104: data <=10'b0000001000; 
      9'd105: data <=10'b0000000100; 
      9'd106: data <=10'b0000001000; 
      9'd107: data <=10'b0000000010; 
      9'd108: data <=10'b0000000001; 
      9'd109: data <=10'b0001000000; 
      9'd110: data <=10'b0000100000; 
      9'd111: data <=10'b0100000000; 
      9'd112: data <=10'b0000000100; 
      9'd113: data <=10'b0000001000; 
      9'd114: data <=10'b0000001000; 
      9'd115: data <=10'b1000000000; 
      9'd116: data <=10'b0000000100; 
      9'd117: data <=10'b0001000000; 
      9'd118: data <=10'b1000000000; 
      9'd119: data <=10'b0000000100; 
      9'd120: data <=10'b0000010000; 
      9'd121: data <=10'b0000100000; 
      9'd122: data <=10'b0001000000; 
      9'd123: data <=10'b0000001000; 
      9'd124: data <=10'b0000001000; 
      9'd125: data <=10'b1000000000; 
      9'd126: data <=10'b0000000100; 
      9'd127: data <=10'b0000001000; 
      9'd128: data <=10'b0001000000; 
      9'd129: data <=10'b0000000001; 
      9'd130: data <=10'b0010000000; 
      9'd131: data <=10'b0100000000; 
      9'd132: data <=10'b0100000000; 
      9'd133: data <=10'b0000010000; 
      9'd134: data <=10'b0000000100; 
      9'd135: data <=10'b0000001000; 
      9'd136: data <=10'b0000010000; 
      9'd137: data <=10'b0000000001; 
      9'd138: data <=10'b0000010000; 
      9'd139: data <=10'b0000000001; 
      9'd140: data <=10'b0000000001; 
      9'd141: data <=10'b0000000001; 
      9'd142: data <=10'b1000000000; 
      9'd143: data <=10'b0000100000; 
      9'd144: data <=10'b1000000000; 
      9'd145: data <=10'b0000100000; 
      9'd146: data <=10'b0000001000; 
      9'd147: data <=10'b0000000010; 
      9'd148: data <=10'b0001000000; 
      9'd149: data <=10'b0000100000; 
      9'd150: data <=10'b0000000010; 
      9'd151: data <=10'b0000000010; 
      9'd152: data <=10'b1000000000; 
      9'd153: data <=10'b0010000000; 
      9'd154: data <=10'b0000000010; 
      9'd155: data <=10'b0010000000; 
      9'd156: data <=10'b0100000000; 
      9'd157: data <=10'b0010000000; 
      9'd158: data <=10'b0000000010; 
      9'd159: data <=10'b0000000001; 
      9'd160: data <=10'b0000000001; 
      9'd161: data <=10'b0000000100; 
      9'd162: data <=10'b0000001000; 
      9'd163: data <=10'b0000001000; 
      9'd164: data <=10'b0000000010; 
      9'd165: data <=10'b0001000000; 
      9'd166: data <=10'b0001000000; 
      9'd167: data <=10'b0000001000; 
      9'd168: data <=10'b0001000000; 
      9'd169: data <=10'b0000001000; 
      9'd170: data <=10'b0100000000; 
      9'd171: data <=10'b0000001000; 
      9'd172: data <=10'b0000010000; 
      9'd173: data <=10'b0000000100; 
      9'd174: data <=10'b1000000000; 
      9'd175: data <=10'b0000001000; 
      9'd176: data <=10'b0000001000; 
      9'd177: data <=10'b0000010000; 
      9'd178: data <=10'b0000100000; 
      9'd179: data <=10'b0000010000; 
      9'd180: data <=10'b0000000100; 
      9'd181: data <=10'b0000001000; 
      9'd182: data <=10'b0000000010; 
      9'd183: data <=10'b0001000000; 
      9'd184: data <=10'b0000000010; 
      9'd185: data <=10'b0001000000; 
      9'd186: data <=10'b0100000000; 
      9'd187: data <=10'b0010000000; 
      9'd188: data <=10'b1000000000; 
      9'd189: data <=10'b0001000000; 
      9'd190: data <=10'b0000000001; 
      9'd191: data <=10'b0100000000; 
      9'd192: data <=10'b0000000100; 
      9'd193: data <=10'b0000000001; 
      9'd194: data <=10'b0000000001; 
      9'd195: data <=10'b0000000010; 
      9'd196: data <=10'b1000000000; 
      9'd197: data <=10'b0000000100; 
      9'd198: data <=10'b1000000000; 
      9'd199: data <=10'b0000000001; 
      9'd200: data <=10'b0000100000; 
      9'd201: data <=10'b0000010000; 
      9'd202: data <=10'b0000001000; 
      9'd203: data <=10'b0010000000; 
      9'd204: data <=10'b0000100000; 
      9'd205: data <=10'b0100000000; 
      9'd206: data <=10'b0010000000; 
      9'd207: data <=10'b0010000000; 
      9'd208: data <=10'b0000010000; 
      9'd209: data <=10'b0000010000; 
      9'd210: data <=10'b0000100000; 
      9'd211: data <=10'b0000000010; 
      9'd212: data <=10'b0001000000; 
      9'd213: data <=10'b0000001000; 
      9'd214: data <=10'b0100000000; 
      9'd215: data <=10'b0010000000; 
      9'd216: data <=10'b0000001000; 
      9'd217: data <=10'b0010000000; 
      9'd218: data <=10'b1000000000; 
      9'd219: data <=10'b0000001000; 
      9'd220: data <=10'b1000000000; 
      9'd221: data <=10'b0010000000; 
      9'd222: data <=10'b0001000000; 
      9'd223: data <=10'b0000000100; 
      9'd224: data <=10'b0000000010; 
      9'd225: data <=10'b0001000000; 
      9'd226: data <=10'b0000100000; 
      9'd227: data <=10'b0000000100; 
      9'd228: data <=10'b0001000000; 
      9'd229: data <=10'b0010000000; 
      9'd230: data <=10'b0000001000; 
      9'd231: data <=10'b0001000000; 
      9'd232: data <=10'b0000010000; 
      9'd233: data <=10'b0100000000; 
      9'd234: data <=10'b1000000000; 
      9'd235: data <=10'b1000000000; 
      9'd236: data <=10'b0100000000; 
      9'd237: data <=10'b0000000010; 
      9'd238: data <=10'b0000001000; 
      9'd239: data <=10'b0010000000; 
      9'd240: data <=10'b0010000000; 
      9'd241: data <=10'b0010000000; 
      9'd242: data <=10'b0000000001; 
      9'd243: data <=10'b0010000000; 
      9'd244: data <=10'b0001000000; 
      9'd245: data <=10'b0000000010; 
      9'd246: data <=10'b0000000001; 
      9'd247: data <=10'b0000100000; 
      9'd248: data <=10'b1000000000; 
      9'd249: data <=10'b0010000000; 
      9'd250: data <=10'b0000001000; 
      9'd251: data <=10'b0010000000; 
      9'd252: data <=10'b1000000000; 
      9'd253: data <=10'b0000100000; 
      9'd254: data <=10'b0000010000; 
      9'd255: data <=10'b0001000000; 
      9'd256: data <=10'b0000000001; 
      9'd257: data <=10'b0000001000; 
      9'd258: data <=10'b0000100000; 
      9'd259: data <=10'b0000100000; 
      9'd260: data <=10'b0000000100; 
      9'd261: data <=10'b0000000100; 
      9'd262: data <=10'b0001000000; 
      9'd263: data <=10'b0000000001; 
      9'd264: data <=10'b0000100000; 
      9'd265: data <=10'b0000000010; 
      9'd266: data <=10'b1000000000; 
      9'd267: data <=10'b0000000010; 
      9'd268: data <=10'b0000000100; 
      9'd269: data <=10'b0000000010; 
      9'd270: data <=10'b0100000000; 
      9'd271: data <=10'b0000010000; 
      9'd272: data <=10'b0000010000; 
      9'd273: data <=10'b0000000100; 
      9'd274: data <=10'b0000001000; 
      9'd275: data <=10'b0000100000; 
      9'd276: data <=10'b0000000010; 
      9'd277: data <=10'b0000100000; 
      9'd278: data <=10'b0000000010; 
      9'd279: data <=10'b0100000000; 
      9'd280: data <=10'b0100000000; 
      9'd281: data <=10'b0100000000; 
      9'd282: data <=10'b0000001000; 
      9'd283: data <=10'b0001000000; 
      9'd284: data <=10'b0000010000; 
      9'd285: data <=10'b0001000000; 
      9'd286: data <=10'b0000000100; 
      9'd287: data <=10'b0100000000; 
      9'd288: data <=10'b0000100000; 
      9'd289: data <=10'b0000001000; 
      9'd290: data <=10'b0000000100; 
      9'd291: data <=10'b0001000000; 
      9'd292: data <=10'b0000010000; 
      9'd293: data <=10'b0001000000; 
      9'd294: data <=10'b0010000000; 
      9'd295: data <=10'b0000100000; 
      9'd296: data <=10'b0010000000; 
      9'd297: data <=10'b0000000100; 
      9'd298: data <=10'b0000010000; 
      9'd299: data <=10'b0000000010; 
      9'd300: data <=10'b0000100000; 
      9'd301: data <=10'b0000000100; 
      9'd302: data <=10'b0000010000; 
      9'd303: data <=10'b0010000000; 
      9'd304: data <=10'b0000100000; 
      9'd305: data <=10'b0000000001; 
      9'd306: data <=10'b0000000100; 
      9'd307: data <=10'b0000100000; 
      9'd308: data <=10'b0000000001; 
      9'd309: data <=10'b1000000000; 
      9'd310: data <=10'b0010000000; 
      9'd311: data <=10'b0000010000; 
      9'd312: data <=10'b0000000001; 
      9'd313: data <=10'b0001000000; 
      9'd314: data <=10'b0100000000; 
      9'd315: data <=10'b1000000000; 
      9'd316: data <=10'b0000001000; 
      9'd317: data <=10'b0000000010; 
      9'd318: data <=10'b0000000100; 
      9'd319: data <=10'b0100000000; 
      9'd320: data <=10'b0100000000; 
      9'd321: data <=10'b0100000000; 
      9'd322: data <=10'b0001000000; 
      9'd323: data <=10'b0000000010; 
      9'd324: data <=10'b0000100000; 
      9'd325: data <=10'b1000000000; 
      9'd326: data <=10'b0000100000; 
      9'd327: data <=10'b0000100000; 
      9'd328: data <=10'b0000001000; 
      9'd329: data <=10'b0100000000; 
      9'd330: data <=10'b0000010000; 
      9'd331: data <=10'b0000001000; 
      9'd332: data <=10'b0000000010; 
      9'd333: data <=10'b0000100000; 
      9'd334: data <=10'b0000010000; 
      9'd335: data <=10'b0000000001; 
      9'd336: data <=10'b0010000000; 
      9'd337: data <=10'b0000000010; 
      9'd338: data <=10'b0100000000; 
      9'd339: data <=10'b0000100000; 
      9'd340: data <=10'b0000100000; 
      9'd341: data <=10'b0001000000; 
      9'd342: data <=10'b0000000010; 
      9'd343: data <=10'b0001000000; 
      9'd344: data <=10'b0001000000; 
      9'd345: data <=10'b1000000000; 
      9'd346: data <=10'b0100000000; 
      9'd347: data <=10'b0010000000; 
      9'd348: data <=10'b0000100000; 
      9'd349: data <=10'b1000000000; 
      9'd350: data <=10'b0000100000; 
      9'd351: data <=10'b0000000010; 
      9'd352: data <=10'b0000010000; 
      9'd353: data <=10'b0000010000; 
      9'd354: data <=10'b0000000010; 
      9'd355: data <=10'b0100000000; 
      9'd356: data <=10'b0000000010; 
      9'd357: data <=10'b0010000000; 
      9'd358: data <=10'b0000010000; 
      9'd359: data <=10'b0000000010; 
      9'd360: data <=10'b0000010000; 
      9'd361: data <=10'b0001000000; 
      9'd362: data <=10'b0000000001; 
      9'd363: data <=10'b0000100000; 
      9'd364: data <=10'b0000001000; 
      9'd365: data <=10'b0010000000; 
      9'd366: data <=10'b0100000000; 
      9'd367: data <=10'b0010000000; 
      9'd368: data <=10'b1000000000; 
      9'd369: data <=10'b0000010000; 
      9'd370: data <=10'b0010000000; 
      9'd371: data <=10'b0010000000; 
      9'd372: data <=10'b0100000000; 
      9'd373: data <=10'b0000100000; 
      9'd374: data <=10'b0000000100; 
      9'd375: data <=10'b0000010000; 
      9'd376: data <=10'b0001000000; 
      9'd377: data <=10'b0001000000; 
      9'd378: data <=10'b0000001000; 
      9'd379: data <=10'b0000100000; 
      9'd380: data <=10'b1000000000; 
      9'd381: data <=10'b0000100000; 
      9'd382: data <=10'b0010000000; 
      9'd383: data <=10'b0010000000; 
      9'd384: data <=10'b0000000100; 
      9'd385: data <=10'b0000000010; 
      9'd386: data <=10'b0000010000; 
      9'd387: data <=10'b0000010000; 
      9'd388: data <=10'b0010000000; 
      9'd389: data <=10'b0000000010; 
      9'd390: data <=10'b0000010000; 
      9'd391: data <=10'b0000100000; 
      9'd392: data <=10'b0000010000; 
      9'd393: data <=10'b0000001000; 
      9'd394: data <=10'b0000000100; 
      9'd395: data <=10'b0010000000; 
      9'd396: data <=10'b0000000001; 
      9'd397: data <=10'b0000010000; 
      9'd398: data <=10'b0100000000; 
      9'd399: data <=10'b0000000010; 
      9'd400: data <=10'b0000000001; 
      9'd401: data <=10'b0000000001; 
      9'd402: data <=10'b0000100000; 
      9'd403: data <=10'b1000000000; 
      9'd404: data <=10'b0000001000; 
      9'd405: data <=10'b0010000000; 
      9'd406: data <=10'b0100000000; 
      9'd407: data <=10'b0000001000; 
      9'd408: data <=10'b0010000000; 
      9'd409: data <=10'b0000000001; 
      9'd410: data <=10'b1000000000; 
      9'd411: data <=10'b0000000010; 
      9'd412: data <=10'b0000010000; 
      9'd413: data <=10'b0000000001; 
      9'd414: data <=10'b0000000010; 
      9'd415: data <=10'b1000000000; 
      9'd416: data <=10'b0010000000; 
      9'd417: data <=10'b1000000000; 
      9'd418: data <=10'b0001000000; 
      9'd419: data <=10'b0000000100; 
      9'd420: data <=10'b0000100000; 
      9'd421: data <=10'b0000010000; 
      9'd422: data <=10'b0001000000; 
      9'd423: data <=10'b0000001000; 
      9'd424: data <=10'b0000000010; 
      9'd425: data <=10'b0000001000; 
      9'd426: data <=10'b0001000000; 
      9'd427: data <=10'b0000000001; 
      9'd428: data <=10'b0000000010; 
      9'd429: data <=10'b0000000001; 
      9'd430: data <=10'b0000010000; 
      9'd431: data <=10'b0000010000; 
      9'd432: data <=10'b0010000000; 
      9'd433: data <=10'b0000000001; 
      9'd434: data <=10'b0000000010; 
      9'd435: data <=10'b0000100000; 
      9'd436: data <=10'b0100000000; 
      9'd437: data <=10'b0000000010; 
      9'd438: data <=10'b0000000100; 
      9'd439: data <=10'b0000000100; 
      9'd440: data <=10'b0000010000; 
      9'd441: data <=10'b0000010000; 
      9'd442: data <=10'b0000010000; 
      9'd443: data <=10'b0001000000; 
      9'd444: data <=10'b1000000000; 
      9'd445: data <=10'b0010000000; 
      9'd446: data <=10'b0000000001; 
      9'd447: data <=10'b0000000001; 
      9'd448: data <=10'b0000000100; 
      9'd449: data <=10'b0100000000; 
      9'd450: data <=10'b0000100000; 
      9'd451: data <=10'b0000000100; 
      9'd452: data <=10'b0000000010; 
      9'd453: data <=10'b0010000000; 
      9'd454: data <=10'b0001000000; 
      9'd455: data <=10'b1000000000; 
      9'd456: data <=10'b0100000000; 
      9'd457: data <=10'b0000000100; 
      9'd458: data <=10'b0100000000; 
      9'd459: data <=10'b0000001000; 
      9'd460: data <=10'b0010000000; 
      9'd461: data <=10'b0010000000; 
      9'd462: data <=10'b0100000000; 
      9'd463: data <=10'b0001000000; 
      9'd464: data <=10'b1000000000; 
      9'd465: data <=10'b0000000010; 
      9'd466: data <=10'b0000000001; 
      9'd467: data <=10'b0010000000; 
      9'd468: data <=10'b0001000000; 
      9'd469: data <=10'b1000000000; 
      9'd470: data <=10'b0000000010; 
      9'd471: data <=10'b1000000000; 
      9'd472: data <=10'b0100000000; 
      9'd473: data <=10'b0001000000; 
      9'd474: data <=10'b0000000100; 
      9'd475: data <=10'b0001000000; 
      9'd476: data <=10'b0000000010; 
      9'd477: data <=10'b0000001000; 
      9'd478: data <=10'b0100000000; 
      9'd479: data <=10'b0000001000; 
      9'd480: data <=10'b0100000000; 
      9'd481: data <=10'b0010000000; 
      9'd482: data <=10'b0000000100; 
      9'd483: data <=10'b0000001000; 
      9'd484: data <=10'b0100000000; 
      9'd485: data <=10'b0000000100; 
      9'd486: data <=10'b0001000000; 
      9'd487: data <=10'b0000000010; 
      9'd488: data <=10'b0000100000; 
      9'd489: data <=10'b0000000100; 
      9'd490: data <=10'b1000000000; 
      9'd491: data <=10'b1000000000; 
      9'd492: data <=10'b0000010000; 
      9'd493: data <=10'b0001000000; 
      default: data<=10'd0;
    endcase 
  end 
endmodule 
