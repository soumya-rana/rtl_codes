`timescale 1ns/1ps 

///////////////////////////////////////////////////////////////////////////////
// Company: Indian Institute of Science, Bengaluru 
// Engineer: Soumya Kanta Rana 
//
// Create Date: 17.11.2021
// Module Name: ROMs for W21 
// Project Name: ELM engine
// Target Devices: xc7a200tfbg484-2
//
////////////////////////////////////////////////////////////////////////////////
module w21_rom8(input [12:0] addr, input clk,  output reg [15:0] data);
  always @ ( posedge clk ) begin 
     case(addr)
      13'd0: data <=16'b1111111110100110; 
      13'd1: data <=16'b1111111110001110; 
      13'd2: data <=16'b0000000010101010; 
      13'd3: data <=16'b0000000001010010; 
      13'd4: data <=16'b1111111110111110; 
      13'd5: data <=16'b1111111111101000; 
      13'd6: data <=16'b1111111111110010; 
      13'd7: data <=16'b0000000000011000; 
      13'd8: data <=16'b0000000001110100; 
      13'd9: data <=16'b1111111111010010; 
      13'd10: data <=16'b1111111101001111; 
      13'd11: data <=16'b0000000001110010; 
      13'd12: data <=16'b1111111101110111; 
      13'd13: data <=16'b0000000000001101; 
      13'd14: data <=16'b0000000010000100; 
      13'd15: data <=16'b1111111101101011; 
      13'd16: data <=16'b1111111111101011; 
      13'd17: data <=16'b0000000001111000; 
      13'd18: data <=16'b1111111110111101; 
      13'd19: data <=16'b0000000010101110; 
      13'd20: data <=16'b0000000010001100; 
      13'd21: data <=16'b1111111110110101; 
      13'd22: data <=16'b0000000000110001; 
      13'd23: data <=16'b0000000000010100; 
      13'd24: data <=16'b1111111111001100; 
      13'd25: data <=16'b1111111110010111; 
      13'd26: data <=16'b1111111111101010; 
      13'd27: data <=16'b0000000011110111; 
      13'd28: data <=16'b1111111110111111; 
      13'd29: data <=16'b1111111111001110; 
      13'd30: data <=16'b0000000000000011; 
      13'd31: data <=16'b1111111101011101; 
      13'd32: data <=16'b0000000000001001; 
      13'd33: data <=16'b1111111110000100; 
      13'd34: data <=16'b1111111111001001; 
      13'd35: data <=16'b0000000010000101; 
      13'd36: data <=16'b0000000001011101; 
      13'd37: data <=16'b0000000000000110; 
      13'd38: data <=16'b0000000001101011; 
      13'd39: data <=16'b0000000011011010; 
      13'd40: data <=16'b1111111110001101; 
      13'd41: data <=16'b0000000001010011; 
      13'd42: data <=16'b0000000001111001; 
      13'd43: data <=16'b0000000001010001; 
      13'd44: data <=16'b0000000001001100; 
      13'd45: data <=16'b0000000001100101; 
      13'd46: data <=16'b0000000000000010; 
      13'd47: data <=16'b0000000001001101; 
      13'd48: data <=16'b0000000010101110; 
      13'd49: data <=16'b0000000001010001; 
      13'd50: data <=16'b1111111111011101; 
      13'd51: data <=16'b0000000001101100; 
      13'd52: data <=16'b0000000001010010; 
      13'd53: data <=16'b1111111111101000; 
      13'd54: data <=16'b1111111111110101; 
      13'd55: data <=16'b0000000010001010; 
      13'd56: data <=16'b0000000011000101; 
      13'd57: data <=16'b0000000001001001; 
      13'd58: data <=16'b0000000011100111; 
      13'd59: data <=16'b0000000001011110; 
      13'd60: data <=16'b0000000000011100; 
      13'd61: data <=16'b1111111101000111; 
      13'd62: data <=16'b1111111101011001; 
      13'd63: data <=16'b0000000000111000; 
      13'd64: data <=16'b0000000001111011; 
      13'd65: data <=16'b0000000000100011; 
      13'd66: data <=16'b0000000000100001; 
      13'd67: data <=16'b0000000001000000; 
      13'd68: data <=16'b0000000001000000; 
      13'd69: data <=16'b0000000001010111; 
      13'd70: data <=16'b1111111111001011; 
      13'd71: data <=16'b1111111111110100; 
      13'd72: data <=16'b0000000001010001; 
      13'd73: data <=16'b0000000000110010; 
      13'd74: data <=16'b1111111111100010; 
      13'd75: data <=16'b0000000000010011; 
      13'd76: data <=16'b1111111111110111; 
      13'd77: data <=16'b0000000000000111; 
      13'd78: data <=16'b0000000000110111; 
      13'd79: data <=16'b1111111101111101; 
      13'd80: data <=16'b1111111101111100; 
      13'd81: data <=16'b1111111101110010; 
      13'd82: data <=16'b1111111110101000; 
      13'd83: data <=16'b1111111111101111; 
      13'd84: data <=16'b0000000001110100; 
      13'd85: data <=16'b0000000011101110; 
      13'd86: data <=16'b1111111111001110; 
      13'd87: data <=16'b0000000000101101; 
      13'd88: data <=16'b0000000001011011; 
      13'd89: data <=16'b0000000000110111; 
      13'd90: data <=16'b0000000010011110; 
      13'd91: data <=16'b1111111111000000; 
      13'd92: data <=16'b1111111111111100; 
      13'd93: data <=16'b1111111100101010; 
      13'd94: data <=16'b0000000001100101; 
      13'd95: data <=16'b1111111111010010; 
      13'd96: data <=16'b1111111110110001; 
      13'd97: data <=16'b0000000000001100; 
      13'd98: data <=16'b1111111110011011; 
      13'd99: data <=16'b0000000000000110; 
      13'd100: data <=16'b0000000001000111; 
      13'd101: data <=16'b0000000010001100; 
      13'd102: data <=16'b0000000000000101; 
      13'd103: data <=16'b1111111110110100; 
      13'd104: data <=16'b0000000000100011; 
      13'd105: data <=16'b0000000010010110; 
      13'd106: data <=16'b0000000001111110; 
      13'd107: data <=16'b0000000010110001; 
      13'd108: data <=16'b0000000010000010; 
      13'd109: data <=16'b1111111111111010; 
      13'd110: data <=16'b1111111111001011; 
      13'd111: data <=16'b0000000000111000; 
      13'd112: data <=16'b1111111111111111; 
      13'd113: data <=16'b1111111110010111; 
      13'd114: data <=16'b1111111111101100; 
      13'd115: data <=16'b1111111111001100; 
      13'd116: data <=16'b0000000000111111; 
      13'd117: data <=16'b1111111110110110; 
      13'd118: data <=16'b0000000010001001; 
      13'd119: data <=16'b1111111110000011; 
      13'd120: data <=16'b0000000001000111; 
      13'd121: data <=16'b0000000010001101; 
      13'd122: data <=16'b1111111111110001; 
      13'd123: data <=16'b0000000000111111; 
      13'd124: data <=16'b1111111111010100; 
      13'd125: data <=16'b1111111111110000; 
      13'd126: data <=16'b0000000001011110; 
      13'd127: data <=16'b1111111110100111; 
      13'd128: data <=16'b1111111111101010; 
      13'd129: data <=16'b0000000010001000; 
      13'd130: data <=16'b1111111111001000; 
      13'd131: data <=16'b0000000011000110; 
      13'd132: data <=16'b0000000000101100; 
      13'd133: data <=16'b1111111111010101; 
      13'd134: data <=16'b1111111011111111; 
      13'd135: data <=16'b0000000010001010; 
      13'd136: data <=16'b1111111101100010; 
      13'd137: data <=16'b1111111100111111; 
      13'd138: data <=16'b1111111111010011; 
      13'd139: data <=16'b0000000000111100; 
      13'd140: data <=16'b0000000001010010; 
      13'd141: data <=16'b0000000001100001; 
      13'd142: data <=16'b0000000001010011; 
      13'd143: data <=16'b1111111111000110; 
      13'd144: data <=16'b0000000001000111; 
      13'd145: data <=16'b0000000000110100; 
      13'd146: data <=16'b0000000000100001; 
      13'd147: data <=16'b0000000000100000; 
      13'd148: data <=16'b1111111110011101; 
      13'd149: data <=16'b1111111111001011; 
      13'd150: data <=16'b1111111101011011; 
      13'd151: data <=16'b0000000000010011; 
      13'd152: data <=16'b0000000001011001; 
      13'd153: data <=16'b1111111100010001; 
      13'd154: data <=16'b1111111100100000; 
      13'd155: data <=16'b0000000000100101; 
      13'd156: data <=16'b1111111101010101; 
      13'd157: data <=16'b0000000000000001; 
      13'd158: data <=16'b0000000001001000; 
      13'd159: data <=16'b1111111111110101; 
      13'd160: data <=16'b1111111111110111; 
      13'd161: data <=16'b0000000001001001; 
      13'd162: data <=16'b0000000001101001; 
      13'd163: data <=16'b1111111111010000; 
      13'd164: data <=16'b0000000000000110; 
      13'd165: data <=16'b1111111110010110; 
      13'd166: data <=16'b1111111101110100; 
      13'd167: data <=16'b1111111101101100; 
      13'd168: data <=16'b0000000000000110; 
      13'd169: data <=16'b1111111110111001; 
      13'd170: data <=16'b1111111101110010; 
      13'd171: data <=16'b1111111111000110; 
      13'd172: data <=16'b1111111101111000; 
      13'd173: data <=16'b0000000000110100; 
      13'd174: data <=16'b0000000001001100; 
      13'd175: data <=16'b0000000010011101; 
      13'd176: data <=16'b0000000000001000; 
      13'd177: data <=16'b1111111111101101; 
      13'd178: data <=16'b1111111111100011; 
      13'd179: data <=16'b1111111110100001; 
      13'd180: data <=16'b0000000001110100; 
      13'd181: data <=16'b0000000000101111; 
      13'd182: data <=16'b1111111111111111; 
      13'd183: data <=16'b0000000000001000; 
      13'd184: data <=16'b1111111110000011; 
      13'd185: data <=16'b1111111110111100; 
      13'd186: data <=16'b0000000001100011; 
      13'd187: data <=16'b1111111110001011; 
      13'd188: data <=16'b0000000001111011; 
      13'd189: data <=16'b0000000010110010; 
      13'd190: data <=16'b1111111111101000; 
      13'd191: data <=16'b0000000001001011; 
      13'd192: data <=16'b1111111111011010; 
      13'd193: data <=16'b0000000000110110; 
      13'd194: data <=16'b0000000000101100; 
      13'd195: data <=16'b1111111111101100; 
      13'd196: data <=16'b1111111111011100; 
      13'd197: data <=16'b1111111101000011; 
      13'd198: data <=16'b1111111110010100; 
      13'd199: data <=16'b1111111111010000; 
      13'd200: data <=16'b0000000000100001; 
      13'd201: data <=16'b1111111110010011; 
      13'd202: data <=16'b1111111110101101; 
      13'd203: data <=16'b0000000010111111; 
      13'd204: data <=16'b1111111111010010; 
      13'd205: data <=16'b1111111110111101; 
      13'd206: data <=16'b1111111110110111; 
      13'd207: data <=16'b1111111110011110; 
      13'd208: data <=16'b0000000001100100; 
      13'd209: data <=16'b0000000000100111; 
      13'd210: data <=16'b0000000000110011; 
      13'd211: data <=16'b0000000000111000; 
      13'd212: data <=16'b0000000010011001; 
      13'd213: data <=16'b1111111110001111; 
      13'd214: data <=16'b1111111110111100; 
      13'd215: data <=16'b0000000001101010; 
      13'd216: data <=16'b0000000000011011; 
      13'd217: data <=16'b0000000001011011; 
      13'd218: data <=16'b0000000001000110; 
      13'd219: data <=16'b0000000000110101; 
      13'd220: data <=16'b0000000000000000; 
      13'd221: data <=16'b1111111111101011; 
      13'd222: data <=16'b0000000000010011; 
      13'd223: data <=16'b0000000001011001; 
      13'd224: data <=16'b0000000001000111; 
      13'd225: data <=16'b0000000001000110; 
      13'd226: data <=16'b0000000000010111; 
      13'd227: data <=16'b1111111111000001; 
      13'd228: data <=16'b0000000001011001; 
      13'd229: data <=16'b0000000010011011; 
      13'd230: data <=16'b0000000000000101; 
      13'd231: data <=16'b0000000000110101; 
      13'd232: data <=16'b0000000000110110; 
      13'd233: data <=16'b1111111110111100; 
      13'd234: data <=16'b0000000001100001; 
      13'd235: data <=16'b1111111111110111; 
      13'd236: data <=16'b1111111110110110; 
      13'd237: data <=16'b1111111111001010; 
      13'd238: data <=16'b0000000000010110; 
      13'd239: data <=16'b0000000001100000; 
      13'd240: data <=16'b1111111110000011; 
      13'd241: data <=16'b1111111111010010; 
      13'd242: data <=16'b0000000001001100; 
      13'd243: data <=16'b0000000000011011; 
      13'd244: data <=16'b1111111111000111; 
      13'd245: data <=16'b1111111111111010; 
      13'd246: data <=16'b0000000010001101; 
      13'd247: data <=16'b1111111101101101; 
      13'd248: data <=16'b1111111111010001; 
      13'd249: data <=16'b0000000000100100; 
      13'd250: data <=16'b1111111110000010; 
      13'd251: data <=16'b1111111111111111; 
      13'd252: data <=16'b1111111111111011; 
      13'd253: data <=16'b1111111110101011; 
      13'd254: data <=16'b1111111110101101; 
      13'd255: data <=16'b0000000000101111; 
      13'd256: data <=16'b0000000000100100; 
      13'd257: data <=16'b0000000000010100; 
      13'd258: data <=16'b1111111110100000; 
      13'd259: data <=16'b1111111111011100; 
      13'd260: data <=16'b1111111110011011; 
      13'd261: data <=16'b0000000000111111; 
      13'd262: data <=16'b1111111111101000; 
      13'd263: data <=16'b0000000010000010; 
      13'd264: data <=16'b1111111111111001; 
      13'd265: data <=16'b0000000001011000; 
      13'd266: data <=16'b1111111100000110; 
      13'd267: data <=16'b0000000000101110; 
      13'd268: data <=16'b1111111110101101; 
      13'd269: data <=16'b1111111101110000; 
      13'd270: data <=16'b0000000000101001; 
      13'd271: data <=16'b1111111110101110; 
      13'd272: data <=16'b0000000000111111; 
      13'd273: data <=16'b1111111111001010; 
      13'd274: data <=16'b0000000000111111; 
      13'd275: data <=16'b0000000011010100; 
      13'd276: data <=16'b1111111101101100; 
      13'd277: data <=16'b1111111111110001; 
      13'd278: data <=16'b0000000010011101; 
      13'd279: data <=16'b0000000001100000; 
      13'd280: data <=16'b0000000000110100; 
      13'd281: data <=16'b1111111110101000; 
      13'd282: data <=16'b1111111111000101; 
      13'd283: data <=16'b1111111101111111; 
      13'd284: data <=16'b1111111110111010; 
      13'd285: data <=16'b0000000001100100; 
      13'd286: data <=16'b0000000001100100; 
      13'd287: data <=16'b0000000000011001; 
      13'd288: data <=16'b1111111111110100; 
      13'd289: data <=16'b1111111110111010; 
      13'd290: data <=16'b0000000010010100; 
      13'd291: data <=16'b0000000000111010; 
      13'd292: data <=16'b1111111101010110; 
      13'd293: data <=16'b0000000001100011; 
      13'd294: data <=16'b1111111111000110; 
      13'd295: data <=16'b1111111111000000; 
      13'd296: data <=16'b0000000000011010; 
      13'd297: data <=16'b0000000000011000; 
      13'd298: data <=16'b0000000010011000; 
      13'd299: data <=16'b1111111101100010; 
      13'd300: data <=16'b1111111111101010; 
      13'd301: data <=16'b0000000000110010; 
      13'd302: data <=16'b1111111111010111; 
      13'd303: data <=16'b1111111110100011; 
      13'd304: data <=16'b0000000000101001; 
      13'd305: data <=16'b0000000001101100; 
      13'd306: data <=16'b1111111101001100; 
      13'd307: data <=16'b1111111110110111; 
      13'd308: data <=16'b1111111111100001; 
      13'd309: data <=16'b0000000000111110; 
      13'd310: data <=16'b1111111110111000; 
      13'd311: data <=16'b1111111011111011; 
      13'd312: data <=16'b1111111111111111; 
      13'd313: data <=16'b1111111110110101; 
      13'd314: data <=16'b0000000000010000; 
      13'd315: data <=16'b0000000000001000; 
      13'd316: data <=16'b1111111101100100; 
      13'd317: data <=16'b0000000000110011; 
      13'd318: data <=16'b0000000000111100; 
      13'd319: data <=16'b0000000000010110; 
      13'd320: data <=16'b1111111111100101; 
      13'd321: data <=16'b0000000000000011; 
      13'd322: data <=16'b1111111110100011; 
      13'd323: data <=16'b1111111111011111; 
      13'd324: data <=16'b0000000000100110; 
      13'd325: data <=16'b0000000010101110; 
      13'd326: data <=16'b0000000000000001; 
      13'd327: data <=16'b1111111111100001; 
      13'd328: data <=16'b0000000010000001; 
      13'd329: data <=16'b0000000010101010; 
      13'd330: data <=16'b0000000001110001; 
      13'd331: data <=16'b0000000001110001; 
      13'd332: data <=16'b0000000000110011; 
      13'd333: data <=16'b0000000000100001; 
      13'd334: data <=16'b1111111111001011; 
      13'd335: data <=16'b0000000010000111; 
      13'd336: data <=16'b1111111111110010; 
      13'd337: data <=16'b1111111111100010; 
      13'd338: data <=16'b0000000001111100; 
      13'd339: data <=16'b0000000001100101; 
      13'd340: data <=16'b1111111110001100; 
      13'd341: data <=16'b0000000010010011; 
      13'd342: data <=16'b0000000000110110; 
      13'd343: data <=16'b0000000010111011; 
      13'd344: data <=16'b0000000000110001; 
      13'd345: data <=16'b0000000000010001; 
      13'd346: data <=16'b0000000000101100; 
      13'd347: data <=16'b1111111111110000; 
      13'd348: data <=16'b0000000000111011; 
      13'd349: data <=16'b1111111110011011; 
      13'd350: data <=16'b1111111101010011; 
      13'd351: data <=16'b0000000000010001; 
      13'd352: data <=16'b0000000001000100; 
      13'd353: data <=16'b0000000001111111; 
      13'd354: data <=16'b0000000000001110; 
      13'd355: data <=16'b0000000001010011; 
      13'd356: data <=16'b0000000000100000; 
      13'd357: data <=16'b0000000001100001; 
      13'd358: data <=16'b0000000001110000; 
      13'd359: data <=16'b1111111110100110; 
      13'd360: data <=16'b1111111110101100; 
      13'd361: data <=16'b0000000000100010; 
      13'd362: data <=16'b0000000000111001; 
      13'd363: data <=16'b0000000001110111; 
      13'd364: data <=16'b1111111110111000; 
      13'd365: data <=16'b1111111111000100; 
      13'd366: data <=16'b1111111101000010; 
      13'd367: data <=16'b1111111111100010; 
      13'd368: data <=16'b1111111111101111; 
      13'd369: data <=16'b1111111110101011; 
      13'd370: data <=16'b0000000000011100; 
      13'd371: data <=16'b0000000000010010; 
      13'd372: data <=16'b1111111111000010; 
      13'd373: data <=16'b0000000001110010; 
      13'd374: data <=16'b1111111100110010; 
      13'd375: data <=16'b1111111111000100; 
      13'd376: data <=16'b0000000000100010; 
      13'd377: data <=16'b1111111111011010; 
      13'd378: data <=16'b1111111111001110; 
      13'd379: data <=16'b1111111111111101; 
      13'd380: data <=16'b0000000001001101; 
      13'd381: data <=16'b0000000001111101; 
      13'd382: data <=16'b0000000000000001; 
      13'd383: data <=16'b0000000000000011; 
      13'd384: data <=16'b0000000001011110; 
      13'd385: data <=16'b0000000000001100; 
      13'd386: data <=16'b0000000001101111; 
      13'd387: data <=16'b0000000000001001; 
      13'd388: data <=16'b1111111111111111; 
      13'd389: data <=16'b1111111111001001; 
      13'd390: data <=16'b0000000001100101; 
      13'd391: data <=16'b0000000011010011; 
      13'd392: data <=16'b1111111111100101; 
      13'd393: data <=16'b1111111111100001; 
      13'd394: data <=16'b1111111101000011; 
      13'd395: data <=16'b0000000000000001; 
      13'd396: data <=16'b0000000010111110; 
      13'd397: data <=16'b1111111111000111; 
      13'd398: data <=16'b1111111110010100; 
      13'd399: data <=16'b1111111111000111; 
      13'd400: data <=16'b1111111110101011; 
      13'd401: data <=16'b0000000001010011; 
      13'd402: data <=16'b1111111110101111; 
      13'd403: data <=16'b1111111111000100; 
      13'd404: data <=16'b0000000000100000; 
      13'd405: data <=16'b0000000001010000; 
      13'd406: data <=16'b0000000000101000; 
      13'd407: data <=16'b0000000010011011; 
      13'd408: data <=16'b0000000000101111; 
      13'd409: data <=16'b1111111110000001; 
      13'd410: data <=16'b1111111111110110; 
      13'd411: data <=16'b0000000000100101; 
      13'd412: data <=16'b1111111110001001; 
      13'd413: data <=16'b1111111111111111; 
      13'd414: data <=16'b1111111111110100; 
      13'd415: data <=16'b0000000010110101; 
      13'd416: data <=16'b0000000010000001; 
      13'd417: data <=16'b0000000000010100; 
      13'd418: data <=16'b1111111111100001; 
      13'd419: data <=16'b0000000000000111; 
      13'd420: data <=16'b0000000000010011; 
      13'd421: data <=16'b1111111111111010; 
      13'd422: data <=16'b1111111111001010; 
      13'd423: data <=16'b1111111110100100; 
      13'd424: data <=16'b0000000000010111; 
      13'd425: data <=16'b0000000001101111; 
      13'd426: data <=16'b1111111111010110; 
      13'd427: data <=16'b1111111101110100; 
      13'd428: data <=16'b1111111110001000; 
      13'd429: data <=16'b1111111111101101; 
      13'd430: data <=16'b1111111111000010; 
      13'd431: data <=16'b0000000011010011; 
      13'd432: data <=16'b0000000011010000; 
      13'd433: data <=16'b0000000000001000; 
      13'd434: data <=16'b1111111110100011; 
      13'd435: data <=16'b0000000000010010; 
      13'd436: data <=16'b1111111111011111; 
      13'd437: data <=16'b1111111111011111; 
      13'd438: data <=16'b1111111110100010; 
      13'd439: data <=16'b1111111110101101; 
      13'd440: data <=16'b1111111111011001; 
      13'd441: data <=16'b1111111101111110; 
      13'd442: data <=16'b0000000001101000; 
      13'd443: data <=16'b0000000001001000; 
      13'd444: data <=16'b0000000001000011; 
      13'd445: data <=16'b0000000001000000; 
      13'd446: data <=16'b0000000000111110; 
      13'd447: data <=16'b0000000000001111; 
      13'd448: data <=16'b0000000001011110; 
      13'd449: data <=16'b0000000000110110; 
      13'd450: data <=16'b0000000010110011; 
      13'd451: data <=16'b1111111111111100; 
      13'd452: data <=16'b0000000010101110; 
      13'd453: data <=16'b0000000000011110; 
      13'd454: data <=16'b1111111111000000; 
      13'd455: data <=16'b1111111111111001; 
      13'd456: data <=16'b1111111111111100; 
      13'd457: data <=16'b0000000001101001; 
      13'd458: data <=16'b0000000001000100; 
      13'd459: data <=16'b1111111101110011; 
      13'd460: data <=16'b1111111110110001; 
      13'd461: data <=16'b1111111111000100; 
      13'd462: data <=16'b1111111111000001; 
      13'd463: data <=16'b1111111110111001; 
      13'd464: data <=16'b0000000000100100; 
      13'd465: data <=16'b0000000001010001; 
      13'd466: data <=16'b1111111111100011; 
      13'd467: data <=16'b0000000000101111; 
      13'd468: data <=16'b0000000010100000; 
      13'd469: data <=16'b1111111110000111; 
      13'd470: data <=16'b0000000000000010; 
      13'd471: data <=16'b0000000000011100; 
      13'd472: data <=16'b1111111110111010; 
      13'd473: data <=16'b0000000000110010; 
      13'd474: data <=16'b0000000001100000; 
      13'd475: data <=16'b1111111110011000; 
      13'd476: data <=16'b1111111110001001; 
      13'd477: data <=16'b1111111111101001; 
      13'd478: data <=16'b0000000001010010; 
      13'd479: data <=16'b0000000000100111; 
      13'd480: data <=16'b0000000010000101; 
      13'd481: data <=16'b1111111111110000; 
      13'd482: data <=16'b0000000010000101; 
      13'd483: data <=16'b1111111110100000; 
      13'd484: data <=16'b0000000000000100; 
      13'd485: data <=16'b1111111101000100; 
      13'd486: data <=16'b0000000001011100; 
      13'd487: data <=16'b1111111111110011; 
      13'd488: data <=16'b0000000000010111; 
      13'd489: data <=16'b0000000010010011; 
      13'd490: data <=16'b0000000000001111; 
      13'd491: data <=16'b0000000001000000; 
      13'd492: data <=16'b1111111111011000; 
      13'd493: data <=16'b0000000000111100; 
      13'd494: data <=16'b1111111110110100; 
      13'd495: data <=16'b1111111110100001; 
      13'd496: data <=16'b1111111110110101; 
      13'd497: data <=16'b1111111111110011; 
      13'd498: data <=16'b1111111110111101; 
      13'd499: data <=16'b1111111111101111; 
      13'd500: data <=16'b0000000001111011; 
      13'd501: data <=16'b0000000001101100; 
      13'd502: data <=16'b0000000011011101; 
      13'd503: data <=16'b0000000001001000; 
      13'd504: data <=16'b1111111110101011; 
      13'd505: data <=16'b1111111101001100; 
      13'd506: data <=16'b1111111110110101; 
      13'd507: data <=16'b1111111110001101; 
      13'd508: data <=16'b0000000000011011; 
      13'd509: data <=16'b0000000001111010; 
      13'd510: data <=16'b0000000000000011; 
      13'd511: data <=16'b1111111110100110; 
      13'd512: data <=16'b1111111110101000; 
      13'd513: data <=16'b0000000010000101; 
      13'd514: data <=16'b1111111111010011; 
      13'd515: data <=16'b1111111110100010; 
      13'd516: data <=16'b0000000001010110; 
      13'd517: data <=16'b0000000010010000; 
      13'd518: data <=16'b0000000000110100; 
      13'd519: data <=16'b1111111110001001; 
      13'd520: data <=16'b0000000001111010; 
      13'd521: data <=16'b1111111111111110; 
      13'd522: data <=16'b1111111111010010; 
      13'd523: data <=16'b1111111111101011; 
      13'd524: data <=16'b1111111111010101; 
      13'd525: data <=16'b1111111110111010; 
      13'd526: data <=16'b1111111101100100; 
      13'd527: data <=16'b1111111110010101; 
      13'd528: data <=16'b0000000000100000; 
      13'd529: data <=16'b0000000000110110; 
      13'd530: data <=16'b1111111100100010; 
      13'd531: data <=16'b0000000001010110; 
      13'd532: data <=16'b0000000000010111; 
      13'd533: data <=16'b0000000001101110; 
      13'd534: data <=16'b1111111011110111; 
      13'd535: data <=16'b0000000000001100; 
      13'd536: data <=16'b0000000010000100; 
      13'd537: data <=16'b0000000010000000; 
      13'd538: data <=16'b0000000001000011; 
      13'd539: data <=16'b0000000001101010; 
      13'd540: data <=16'b1111111100111010; 
      13'd541: data <=16'b1111111101111001; 
      13'd542: data <=16'b0000000010011101; 
      13'd543: data <=16'b0000000000010000; 
      13'd544: data <=16'b1111111110000001; 
      13'd545: data <=16'b1111111111110000; 
      13'd546: data <=16'b1111111110110110; 
      13'd547: data <=16'b1111111111111001; 
      13'd548: data <=16'b0000000001010111; 
      13'd549: data <=16'b0000000001010101; 
      13'd550: data <=16'b1111111110001001; 
      13'd551: data <=16'b0000000010011010; 
      13'd552: data <=16'b0000000001001110; 
      13'd553: data <=16'b1111111110100010; 
      13'd554: data <=16'b1111111111001100; 
      13'd555: data <=16'b1111111110111000; 
      13'd556: data <=16'b1111111111100011; 
      13'd557: data <=16'b0000000001100110; 
      13'd558: data <=16'b0000000001010100; 
      13'd559: data <=16'b1111111111001010; 
      13'd560: data <=16'b0000000001001000; 
      13'd561: data <=16'b1111111111111100; 
      13'd562: data <=16'b0000000000010001; 
      13'd563: data <=16'b1111111111010011; 
      13'd564: data <=16'b0000000000010001; 
      13'd565: data <=16'b1111111110011111; 
      13'd566: data <=16'b1111111111011100; 
      13'd567: data <=16'b1111111111100101; 
      13'd568: data <=16'b1111111110010110; 
      13'd569: data <=16'b0000000001010100; 
      13'd570: data <=16'b0000000001000100; 
      13'd571: data <=16'b0000000010011101; 
      13'd572: data <=16'b0000000010001101; 
      13'd573: data <=16'b1111111111010001; 
      13'd574: data <=16'b1111111101100100; 
      13'd575: data <=16'b1111111111010011; 
      13'd576: data <=16'b1111111111110010; 
      13'd577: data <=16'b0000000010001010; 
      13'd578: data <=16'b1111111111000001; 
      13'd579: data <=16'b0000000000110001; 
      13'd580: data <=16'b1111111111000101; 
      13'd581: data <=16'b1111111111110111; 
      13'd582: data <=16'b0000000000100001; 
      13'd583: data <=16'b0000000000111010; 
      13'd584: data <=16'b0000000001011010; 
      13'd585: data <=16'b0000000000111101; 
      13'd586: data <=16'b0000000001010111; 
      13'd587: data <=16'b0000000000101101; 
      13'd588: data <=16'b1111111111111100; 
      13'd589: data <=16'b1111111101101110; 
      13'd590: data <=16'b1111111101101010; 
      13'd591: data <=16'b1111111111111010; 
      13'd592: data <=16'b1111111110110110; 
      13'd593: data <=16'b1111111110111110; 
      13'd594: data <=16'b1111111111011100; 
      13'd595: data <=16'b1111111110111011; 
      13'd596: data <=16'b1111111110011001; 
      13'd597: data <=16'b0000000001000011; 
      13'd598: data <=16'b0000000001100101; 
      13'd599: data <=16'b1111111111010000; 
      13'd600: data <=16'b0000000001010101; 
      13'd601: data <=16'b0000000000010010; 
      13'd602: data <=16'b0000000010101101; 
      13'd603: data <=16'b0000000000001100; 
      13'd604: data <=16'b1111111111101110; 
      13'd605: data <=16'b1111111110111100; 
      13'd606: data <=16'b0000000000010101; 
      13'd607: data <=16'b0000000000000010; 
      13'd608: data <=16'b0000000001101001; 
      13'd609: data <=16'b1111111110001111; 
      13'd610: data <=16'b0000000000110110; 
      13'd611: data <=16'b0000000000101000; 
      13'd612: data <=16'b0000000001001011; 
      13'd613: data <=16'b0000000000110000; 
      13'd614: data <=16'b0000000000100001; 
      13'd615: data <=16'b0000000000011111; 
      13'd616: data <=16'b0000000001000111; 
      13'd617: data <=16'b0000000001110100; 
      13'd618: data <=16'b0000000001011011; 
      13'd619: data <=16'b0000000010101001; 
      13'd620: data <=16'b1111111111000101; 
      13'd621: data <=16'b0000000000001101; 
      13'd622: data <=16'b1111111111000001; 
      13'd623: data <=16'b0000000001110010; 
      13'd624: data <=16'b1111111111100000; 
      13'd625: data <=16'b0000000000011101; 
      13'd626: data <=16'b1111111111100001; 
      13'd627: data <=16'b0000000010010010; 
      13'd628: data <=16'b1111111110100001; 
      13'd629: data <=16'b1111111110100111; 
      13'd630: data <=16'b1111111111000110; 
      13'd631: data <=16'b1111111111101101; 
      13'd632: data <=16'b0000000010010000; 
      13'd633: data <=16'b0000000000011111; 
      13'd634: data <=16'b1111111111011111; 
      13'd635: data <=16'b0000000000100101; 
      13'd636: data <=16'b1111111111101011; 
      13'd637: data <=16'b0000000000001111; 
      13'd638: data <=16'b0000000000111111; 
      13'd639: data <=16'b1111111111101110; 
      13'd640: data <=16'b1111111101100011; 
      13'd641: data <=16'b0000000001000011; 
      13'd642: data <=16'b1111111101011100; 
      13'd643: data <=16'b1111111110110111; 
      13'd644: data <=16'b1111111111011011; 
      13'd645: data <=16'b0000000001110111; 
      13'd646: data <=16'b0000000010010101; 
      13'd647: data <=16'b1111111111011111; 
      13'd648: data <=16'b1111111110100010; 
      13'd649: data <=16'b1111111111001100; 
      13'd650: data <=16'b1111111100101011; 
      13'd651: data <=16'b1111111111001010; 
      13'd652: data <=16'b0000000001010110; 
      13'd653: data <=16'b1111111101001011; 
      13'd654: data <=16'b1111111110101010; 
      13'd655: data <=16'b1111111110010001; 
      13'd656: data <=16'b1111111110111010; 
      13'd657: data <=16'b0000000000000010; 
      13'd658: data <=16'b0000000000100100; 
      13'd659: data <=16'b0000000000101010; 
      13'd660: data <=16'b0000000000111110; 
      13'd661: data <=16'b1111111101101100; 
      13'd662: data <=16'b1111111110101001; 
      13'd663: data <=16'b1111111111101100; 
      13'd664: data <=16'b0000000000011001; 
      13'd665: data <=16'b1111111111001011; 
      13'd666: data <=16'b1111111110010100; 
      13'd667: data <=16'b1111111111000110; 
      13'd668: data <=16'b1111111101111000; 
      13'd669: data <=16'b0000000000011011; 
      13'd670: data <=16'b1111111111011111; 
      13'd671: data <=16'b0000000000101000; 
      13'd672: data <=16'b0000000001010110; 
      13'd673: data <=16'b1111111101100000; 
      13'd674: data <=16'b1111111111000111; 
      13'd675: data <=16'b0000000011000101; 
      13'd676: data <=16'b0000000000100000; 
      13'd677: data <=16'b1111111111001101; 
      13'd678: data <=16'b1111111111010000; 
      13'd679: data <=16'b1111111110110110; 
      13'd680: data <=16'b1111111111001010; 
      13'd681: data <=16'b0000000000001110; 
      13'd682: data <=16'b1111111110011001; 
      13'd683: data <=16'b0000000000111001; 
      13'd684: data <=16'b0000000001100011; 
      13'd685: data <=16'b1111111110110101; 
      13'd686: data <=16'b1111111111101000; 
      13'd687: data <=16'b0000000001100110; 
      13'd688: data <=16'b1111111111100111; 
      13'd689: data <=16'b0000000001010001; 
      13'd690: data <=16'b1111111101110101; 
      13'd691: data <=16'b0000000000000101; 
      13'd692: data <=16'b0000000000000110; 
      13'd693: data <=16'b0000000001100011; 
      13'd694: data <=16'b0000000000100110; 
      13'd695: data <=16'b0000000000001110; 
      13'd696: data <=16'b0000000000010110; 
      13'd697: data <=16'b1111111111011111; 
      13'd698: data <=16'b0000000001011000; 
      13'd699: data <=16'b0000000001100111; 
      13'd700: data <=16'b0000000000000110; 
      13'd701: data <=16'b0000000010010100; 
      13'd702: data <=16'b1111111110110110; 
      13'd703: data <=16'b1111111111011101; 
      13'd704: data <=16'b0000000001001110; 
      13'd705: data <=16'b1111111111000011; 
      13'd706: data <=16'b1111111111110000; 
      13'd707: data <=16'b0000000010111101; 
      13'd708: data <=16'b0000000010111001; 
      13'd709: data <=16'b1111111111011001; 
      13'd710: data <=16'b0000000000010001; 
      13'd711: data <=16'b0000000001011101; 
      13'd712: data <=16'b1111111110100111; 
      13'd713: data <=16'b0000000000100011; 
      13'd714: data <=16'b0000000010011010; 
      13'd715: data <=16'b1111111110101110; 
      13'd716: data <=16'b1111111111111000; 
      13'd717: data <=16'b1111111110101001; 
      13'd718: data <=16'b1111111111110001; 
      13'd719: data <=16'b0000000001110000; 
      13'd720: data <=16'b0000000010101001; 
      13'd721: data <=16'b0000000000111011; 
      13'd722: data <=16'b1111111110000110; 
      13'd723: data <=16'b1111111110110111; 
      13'd724: data <=16'b0000000000001110; 
      13'd725: data <=16'b1111111101110001; 
      13'd726: data <=16'b1111111101110010; 
      13'd727: data <=16'b0000000000011000; 
      13'd728: data <=16'b1111111111100001; 
      13'd729: data <=16'b1111111111101110; 
      13'd730: data <=16'b1111111110001110; 
      13'd731: data <=16'b1111111111011111; 
      13'd732: data <=16'b1111111111001000; 
      13'd733: data <=16'b1111111111111011; 
      13'd734: data <=16'b0000000010010100; 
      13'd735: data <=16'b1111111110101110; 
      13'd736: data <=16'b1111111111110110; 
      13'd737: data <=16'b1111111111101000; 
      13'd738: data <=16'b1111111110100001; 
      13'd739: data <=16'b0000000001010010; 
      13'd740: data <=16'b0000000001111101; 
      13'd741: data <=16'b0000000000111000; 
      13'd742: data <=16'b0000000000111001; 
      13'd743: data <=16'b0000000000010111; 
      13'd744: data <=16'b1111111111101010; 
      13'd745: data <=16'b1111111111110111; 
      13'd746: data <=16'b1111111110010110; 
      13'd747: data <=16'b0000000001001001; 
      13'd748: data <=16'b0000000011000101; 
      13'd749: data <=16'b1111111111010001; 
      13'd750: data <=16'b0000000001000010; 
      13'd751: data <=16'b1111111110100111; 
      13'd752: data <=16'b0000000000011001; 
      13'd753: data <=16'b1111111110111001; 
      13'd754: data <=16'b0000000001101011; 
      13'd755: data <=16'b1111111111101100; 
      13'd756: data <=16'b0000000000011110; 
      13'd757: data <=16'b0000000001101000; 
      13'd758: data <=16'b0000000001011011; 
      13'd759: data <=16'b0000000000110010; 
      13'd760: data <=16'b0000000001100111; 
      13'd761: data <=16'b1111111111001010; 
      13'd762: data <=16'b0000000000001101; 
      13'd763: data <=16'b1111111101010011; 
      13'd764: data <=16'b0000000000111001; 
      13'd765: data <=16'b0000000000110111; 
      13'd766: data <=16'b0000000001011110; 
      13'd767: data <=16'b1111111111111000; 
      13'd768: data <=16'b1111111111011010; 
      13'd769: data <=16'b1111111110101110; 
      13'd770: data <=16'b1111111101101011; 
      13'd771: data <=16'b1111111110010010; 
      13'd772: data <=16'b0000000001010010; 
      13'd773: data <=16'b1111111101100100; 
      13'd774: data <=16'b1111111111011000; 
      13'd775: data <=16'b1111111111100011; 
      13'd776: data <=16'b1111111111010001; 
      13'd777: data <=16'b0000000010000010; 
      13'd778: data <=16'b0000000001010001; 
      13'd779: data <=16'b1111111110001100; 
      13'd780: data <=16'b1111111101100101; 
      13'd781: data <=16'b1111111111101110; 
      13'd782: data <=16'b0000000001110010; 
      13'd783: data <=16'b1111111111111010; 
      13'd784: data <=16'b1111111111001010; 
      13'd785: data <=16'b1111111101110011; 
      13'd786: data <=16'b0000000000100000; 
      13'd787: data <=16'b1111111111100110; 
      13'd788: data <=16'b0000000001111110; 
      13'd789: data <=16'b0000000000111011; 
      13'd790: data <=16'b1111111100111110; 
      13'd791: data <=16'b0000000001000101; 
      13'd792: data <=16'b1111111111011100; 
      13'd793: data <=16'b0000000001010100; 
      13'd794: data <=16'b0000000001001000; 
      13'd795: data <=16'b1111111111010000; 
      13'd796: data <=16'b1111111110111110; 
      13'd797: data <=16'b1111111100111101; 
      13'd798: data <=16'b0000000001001110; 
      13'd799: data <=16'b1111111111110100; 
      13'd800: data <=16'b0000000000010010; 
      13'd801: data <=16'b1111111110011000; 
      13'd802: data <=16'b0000000000000111; 
      13'd803: data <=16'b0000000001010010; 
      13'd804: data <=16'b0000000000011100; 
      13'd805: data <=16'b0000000000000110; 
      13'd806: data <=16'b1111111101110010; 
      13'd807: data <=16'b1111111110101111; 
      13'd808: data <=16'b0000000001010100; 
      13'd809: data <=16'b0000000001001011; 
      13'd810: data <=16'b1111111111110101; 
      13'd811: data <=16'b1111111100010010; 
      13'd812: data <=16'b0000000000110110; 
      13'd813: data <=16'b1111111110110011; 
      13'd814: data <=16'b1111111110010010; 
      13'd815: data <=16'b1111111101110110; 
      13'd816: data <=16'b0000000000101110; 
      13'd817: data <=16'b1111111111000000; 
      13'd818: data <=16'b1111111110100011; 
      13'd819: data <=16'b1111111111001011; 
      13'd820: data <=16'b1111111110110011; 
      13'd821: data <=16'b0000000001110011; 
      13'd822: data <=16'b1111111111000011; 
      13'd823: data <=16'b1111111110110110; 
      13'd824: data <=16'b1111111110011001; 
      13'd825: data <=16'b1111111111001110; 
      13'd826: data <=16'b1111111111011111; 
      13'd827: data <=16'b0000000001111101; 
      13'd828: data <=16'b0000000001011001; 
      13'd829: data <=16'b1111111111111101; 
      13'd830: data <=16'b0000000001111001; 
      13'd831: data <=16'b1111111111000001; 
      13'd832: data <=16'b1111111111100110; 
      13'd833: data <=16'b0000000001001010; 
      13'd834: data <=16'b0000000000000111; 
      13'd835: data <=16'b0000000000101011; 
      13'd836: data <=16'b1111111111101011; 
      13'd837: data <=16'b1111111100110000; 
      13'd838: data <=16'b1111111110111001; 
      13'd839: data <=16'b1111111111111011; 
      13'd840: data <=16'b0000000000001100; 
      13'd841: data <=16'b1111111110100011; 
      13'd842: data <=16'b0000000000101011; 
      13'd843: data <=16'b0000000001001100; 
      13'd844: data <=16'b1111111101101011; 
      13'd845: data <=16'b0000000001001111; 
      13'd846: data <=16'b0000000010011111; 
      13'd847: data <=16'b0000000000001100; 
      13'd848: data <=16'b1111111101001110; 
      13'd849: data <=16'b1111111110111110; 
      13'd850: data <=16'b1111111110110000; 
      13'd851: data <=16'b0000000000101101; 
      13'd852: data <=16'b1111111111010011; 
      13'd853: data <=16'b0000000001011101; 
      13'd854: data <=16'b0000000001101100; 
      13'd855: data <=16'b0000000000111001; 
      13'd856: data <=16'b1111111111100011; 
      13'd857: data <=16'b0000000010110101; 
      13'd858: data <=16'b1111111110100111; 
      13'd859: data <=16'b0000000000110110; 
      13'd860: data <=16'b1111111110011011; 
      13'd861: data <=16'b0000000000010001; 
      13'd862: data <=16'b1111111111111101; 
      13'd863: data <=16'b0000000000001110; 
      13'd864: data <=16'b0000000010010111; 
      13'd865: data <=16'b0000000000110110; 
      13'd866: data <=16'b0000000000110001; 
      13'd867: data <=16'b0000000000010001; 
      13'd868: data <=16'b0000000001100111; 
      13'd869: data <=16'b1111111111110001; 
      13'd870: data <=16'b0000000001101011; 
      13'd871: data <=16'b0000000000100011; 
      13'd872: data <=16'b1111111101000010; 
      13'd873: data <=16'b0000000010001010; 
      13'd874: data <=16'b1111111111001010; 
      13'd875: data <=16'b0000000010110010; 
      13'd876: data <=16'b1111111111011100; 
      13'd877: data <=16'b1111111111001101; 
      13'd878: data <=16'b1111111110011111; 
      13'd879: data <=16'b1111111110101111; 
      13'd880: data <=16'b0000000000111000; 
      13'd881: data <=16'b0000000000101110; 
      13'd882: data <=16'b0000000001101000; 
      13'd883: data <=16'b1111111111101111; 
      13'd884: data <=16'b1111111101010000; 
      13'd885: data <=16'b1111111111111011; 
      13'd886: data <=16'b1111111111101111; 
      13'd887: data <=16'b1111111111001001; 
      13'd888: data <=16'b1111111100010001; 
      13'd889: data <=16'b1111111111011010; 
      13'd890: data <=16'b1111111111110100; 
      13'd891: data <=16'b1111111110101111; 
      13'd892: data <=16'b0000000001011111; 
      13'd893: data <=16'b1111111111001111; 
      13'd894: data <=16'b0000000000001111; 
      13'd895: data <=16'b0000000000011000; 
      13'd896: data <=16'b1111111110000111; 
      13'd897: data <=16'b1111111110101001; 
      13'd898: data <=16'b0000000001110010; 
      13'd899: data <=16'b1111111100101100; 
      13'd900: data <=16'b1111111111001000; 
      13'd901: data <=16'b1111111111101100; 
      13'd902: data <=16'b0000000000001101; 
      13'd903: data <=16'b1111111111111010; 
      13'd904: data <=16'b0000000000100110; 
      13'd905: data <=16'b0000000000001100; 
      13'd906: data <=16'b1111111111010001; 
      13'd907: data <=16'b0000000001011101; 
      13'd908: data <=16'b0000000001011000; 
      13'd909: data <=16'b0000000001011100; 
      13'd910: data <=16'b1111111110101110; 
      13'd911: data <=16'b1111111110000010; 
      13'd912: data <=16'b0000000010100111; 
      13'd913: data <=16'b0000000000111001; 
      13'd914: data <=16'b0000000010010110; 
      13'd915: data <=16'b1111111101101011; 
      13'd916: data <=16'b1111111111001111; 
      13'd917: data <=16'b0000000000111100; 
      13'd918: data <=16'b0000000000101111; 
      13'd919: data <=16'b1111111110101100; 
      13'd920: data <=16'b1111111110110011; 
      13'd921: data <=16'b1111111111100001; 
      13'd922: data <=16'b1111111111101010; 
      13'd923: data <=16'b1111111101111100; 
      13'd924: data <=16'b1111111111101101; 
      13'd925: data <=16'b1111111110000100; 
      13'd926: data <=16'b1111111111010011; 
      13'd927: data <=16'b1111111111011011; 
      13'd928: data <=16'b1111111111010011; 
      13'd929: data <=16'b0000000010001011; 
      13'd930: data <=16'b1111111111001000; 
      13'd931: data <=16'b1111111111001101; 
      13'd932: data <=16'b0000000001011110; 
      13'd933: data <=16'b1111111100100001; 
      13'd934: data <=16'b1111111111101011; 
      13'd935: data <=16'b0000000011100110; 
      13'd936: data <=16'b1111111111000000; 
      13'd937: data <=16'b0000000001000110; 
      13'd938: data <=16'b0000000000010111; 
      13'd939: data <=16'b0000000000010101; 
      13'd940: data <=16'b1111111110101010; 
      13'd941: data <=16'b1111111111011100; 
      13'd942: data <=16'b0000000000111100; 
      13'd943: data <=16'b1111111111111111; 
      13'd944: data <=16'b0000000010010111; 
      13'd945: data <=16'b1111111111001000; 
      13'd946: data <=16'b0000000001000000; 
      13'd947: data <=16'b1111111110010000; 
      13'd948: data <=16'b1111111111111011; 
      13'd949: data <=16'b0000000001111001; 
      13'd950: data <=16'b0000000000000010; 
      13'd951: data <=16'b0000000000100111; 
      13'd952: data <=16'b1111111111111001; 
      13'd953: data <=16'b1111111111001110; 
      13'd954: data <=16'b1111111111101001; 
      13'd955: data <=16'b1111111110110101; 
      13'd956: data <=16'b1111111111110011; 
      13'd957: data <=16'b1111111110111100; 
      13'd958: data <=16'b0000000000101011; 
      13'd959: data <=16'b1111111110011010; 
      13'd960: data <=16'b1111111111011100; 
      13'd961: data <=16'b1111111111000111; 
      13'd962: data <=16'b0000000001010100; 
      13'd963: data <=16'b0000000001011001; 
      13'd964: data <=16'b1111111110001100; 
      13'd965: data <=16'b0000000001101011; 
      13'd966: data <=16'b1111111111111000; 
      13'd967: data <=16'b0000000000001010; 
      13'd968: data <=16'b1111111111101011; 
      13'd969: data <=16'b1111111101001000; 
      13'd970: data <=16'b1111111101101101; 
      13'd971: data <=16'b0000000000011010; 
      13'd972: data <=16'b1111111110110000; 
      13'd973: data <=16'b1111111111111000; 
      13'd974: data <=16'b0000000001000001; 
      13'd975: data <=16'b0000000001100110; 
      13'd976: data <=16'b0000000001111001; 
      13'd977: data <=16'b1111111111101010; 
      13'd978: data <=16'b0000000001101001; 
      13'd979: data <=16'b1111111100110101; 
      13'd980: data <=16'b0000000011000011; 
      13'd981: data <=16'b0000000001100110; 
      13'd982: data <=16'b0000000000011010; 
      13'd983: data <=16'b0000000001011011; 
      13'd984: data <=16'b0000000000001110; 
      13'd985: data <=16'b0000000000011100; 
      13'd986: data <=16'b1111111111101110; 
      13'd987: data <=16'b1111111110100101; 
      13'd988: data <=16'b0000000010000100; 
      13'd989: data <=16'b1111111111001011; 
      13'd990: data <=16'b1111111111011100; 
      13'd991: data <=16'b0000000001011000; 
      13'd992: data <=16'b0000000000001010; 
      13'd993: data <=16'b0000000000100110; 
      13'd994: data <=16'b0000000000011010; 
      13'd995: data <=16'b0000000000011110; 
      13'd996: data <=16'b0000000001111110; 
      13'd997: data <=16'b1111111111000101; 
      13'd998: data <=16'b1111111110111010; 
      13'd999: data <=16'b1111111101101100; 
      13'd1000: data <=16'b0000000010111101; 
      13'd1001: data <=16'b0000000001000010; 
      13'd1002: data <=16'b1111111111101111; 
      13'd1003: data <=16'b1111111111101000; 
      13'd1004: data <=16'b1111111110111111; 
      13'd1005: data <=16'b1111111110101101; 
      13'd1006: data <=16'b0000000001011010; 
      13'd1007: data <=16'b1111111110100110; 
      13'd1008: data <=16'b1111111110111101; 
      13'd1009: data <=16'b1111111110011111; 
      13'd1010: data <=16'b1111111111000011; 
      13'd1011: data <=16'b1111111111010011; 
      13'd1012: data <=16'b1111111110010011; 
      13'd1013: data <=16'b1111111110111101; 
      13'd1014: data <=16'b1111111111100100; 
      13'd1015: data <=16'b1111111110111111; 
      13'd1016: data <=16'b0000000000000101; 
      13'd1017: data <=16'b1111111111011111; 
      13'd1018: data <=16'b1111111111101111; 
      13'd1019: data <=16'b1111111111000111; 
      13'd1020: data <=16'b1111111111111101; 
      13'd1021: data <=16'b0000000001001010; 
      13'd1022: data <=16'b1111111111101001; 
      13'd1023: data <=16'b1111111110001001; 
      13'd1024: data <=16'b1111111110000000; 
      13'd1025: data <=16'b1111111111000110; 
      13'd1026: data <=16'b1111111111100010; 
      13'd1027: data <=16'b0000000001011001; 
      13'd1028: data <=16'b1111111111000110; 
      13'd1029: data <=16'b1111111111110100; 
      13'd1030: data <=16'b0000000001101110; 
      13'd1031: data <=16'b1111111110101101; 
      13'd1032: data <=16'b0000000010101000; 
      13'd1033: data <=16'b0000000000001100; 
      13'd1034: data <=16'b1111111110111101; 
      13'd1035: data <=16'b0000000001111101; 
      13'd1036: data <=16'b1111111111000011; 
      13'd1037: data <=16'b1111111111100101; 
      13'd1038: data <=16'b0000000000001000; 
      13'd1039: data <=16'b0000000001111001; 
      13'd1040: data <=16'b0000000010000010; 
      13'd1041: data <=16'b1111111111101001; 
      13'd1042: data <=16'b0000000010100000; 
      13'd1043: data <=16'b0000000001101000; 
      13'd1044: data <=16'b0000000001011010; 
      13'd1045: data <=16'b1111111110010001; 
      13'd1046: data <=16'b0000000000001101; 
      13'd1047: data <=16'b0000000001000110; 
      13'd1048: data <=16'b1111111111011000; 
      13'd1049: data <=16'b1111111110010110; 
      13'd1050: data <=16'b1111111111111110; 
      13'd1051: data <=16'b1111111110011000; 
      13'd1052: data <=16'b1111111110101011; 
      13'd1053: data <=16'b1111111110001111; 
      13'd1054: data <=16'b1111111101011111; 
      13'd1055: data <=16'b0000000000101001; 
      13'd1056: data <=16'b1111111110010010; 
      13'd1057: data <=16'b1111111110010100; 
      13'd1058: data <=16'b0000000000100111; 
      13'd1059: data <=16'b1111111110101101; 
      13'd1060: data <=16'b1111111100110100; 
      13'd1061: data <=16'b1111111100100111; 
      13'd1062: data <=16'b0000000001010010; 
      13'd1063: data <=16'b1111111111011110; 
      13'd1064: data <=16'b1111111111011110; 
      13'd1065: data <=16'b0000000000010001; 
      13'd1066: data <=16'b1111111110010101; 
      13'd1067: data <=16'b1111111101111111; 
      13'd1068: data <=16'b1111111101100110; 
      13'd1069: data <=16'b0000000000110101; 
      13'd1070: data <=16'b0000000001001101; 
      13'd1071: data <=16'b0000000001000100; 
      13'd1072: data <=16'b0000000000111000; 
      13'd1073: data <=16'b0000000000000100; 
      13'd1074: data <=16'b1111111110101101; 
      13'd1075: data <=16'b0000000011000010; 
      13'd1076: data <=16'b0000000001110000; 
      13'd1077: data <=16'b0000000000000111; 
      13'd1078: data <=16'b1111111100110100; 
      13'd1079: data <=16'b0000000000101100; 
      13'd1080: data <=16'b1111111111111111; 
      13'd1081: data <=16'b0000000000111110; 
      13'd1082: data <=16'b0000000010010101; 
      13'd1083: data <=16'b0000000001100011; 
      13'd1084: data <=16'b0000000010001010; 
      13'd1085: data <=16'b1111111110110000; 
      13'd1086: data <=16'b0000000000010100; 
      13'd1087: data <=16'b0000000011001110; 
      13'd1088: data <=16'b1111111101010110; 
      13'd1089: data <=16'b1111111110101100; 
      13'd1090: data <=16'b1111111111101001; 
      13'd1091: data <=16'b1111111110101100; 
      13'd1092: data <=16'b0000000000001111; 
      13'd1093: data <=16'b0000000001111011; 
      13'd1094: data <=16'b0000000010001001; 
      13'd1095: data <=16'b0000000000000010; 
      13'd1096: data <=16'b0000000001100101; 
      13'd1097: data <=16'b0000000010110101; 
      13'd1098: data <=16'b0000000001000010; 
      13'd1099: data <=16'b1111111100011011; 
      13'd1100: data <=16'b1111111111011000; 
      13'd1101: data <=16'b1111111111110100; 
      13'd1102: data <=16'b1111111110111110; 
      13'd1103: data <=16'b1111111110000000; 
      13'd1104: data <=16'b1111111111001110; 
      13'd1105: data <=16'b0000000000010111; 
      13'd1106: data <=16'b1111111111110101; 
      13'd1107: data <=16'b1111111101110101; 
      13'd1108: data <=16'b1111111111001000; 
      13'd1109: data <=16'b0000000010000100; 
      13'd1110: data <=16'b0000000001101101; 
      13'd1111: data <=16'b1111111110111100; 
      13'd1112: data <=16'b0000000010011001; 
      13'd1113: data <=16'b1111111111010110; 
      13'd1114: data <=16'b0000000010000110; 
      13'd1115: data <=16'b0000000011011110; 
      13'd1116: data <=16'b1111111111010101; 
      13'd1117: data <=16'b0000000000011000; 
      13'd1118: data <=16'b0000000001011101; 
      13'd1119: data <=16'b0000000001001000; 
      13'd1120: data <=16'b0000000001111110; 
      13'd1121: data <=16'b0000000000010110; 
      13'd1122: data <=16'b1111111110111000; 
      13'd1123: data <=16'b0000000000100110; 
      13'd1124: data <=16'b1111111111110000; 
      13'd1125: data <=16'b0000000000011011; 
      13'd1126: data <=16'b1111111110001010; 
      13'd1127: data <=16'b0000000001001100; 
      13'd1128: data <=16'b1111111101001111; 
      13'd1129: data <=16'b1111111111110101; 
      13'd1130: data <=16'b0000000000001100; 
      13'd1131: data <=16'b0000000000011101; 
      13'd1132: data <=16'b0000000000011010; 
      13'd1133: data <=16'b0000000000111101; 
      13'd1134: data <=16'b1111111110100111; 
      13'd1135: data <=16'b1111111111111101; 
      13'd1136: data <=16'b0000000010101101; 
      13'd1137: data <=16'b1111111111011001; 
      13'd1138: data <=16'b1111111111101101; 
      13'd1139: data <=16'b1111111111111100; 
      13'd1140: data <=16'b0000000000011000; 
      13'd1141: data <=16'b0000000000001011; 
      13'd1142: data <=16'b1111111111100110; 
      13'd1143: data <=16'b1111111110111010; 
      13'd1144: data <=16'b0000000001000101; 
      13'd1145: data <=16'b0000000001000100; 
      13'd1146: data <=16'b1111111110101000; 
      13'd1147: data <=16'b0000000001110111; 
      13'd1148: data <=16'b0000000000111101; 
      13'd1149: data <=16'b1111111110100100; 
      13'd1150: data <=16'b0000000000101111; 
      13'd1151: data <=16'b1111111110101101; 
      13'd1152: data <=16'b0000000000001100; 
      13'd1153: data <=16'b1111111111110000; 
      13'd1154: data <=16'b1111111111110001; 
      13'd1155: data <=16'b0000000001000001; 
      13'd1156: data <=16'b0000000000101101; 
      13'd1157: data <=16'b0000000001101001; 
      13'd1158: data <=16'b0000000000111110; 
      13'd1159: data <=16'b0000000000010000; 
      13'd1160: data <=16'b0000000000000010; 
      13'd1161: data <=16'b0000000001001001; 
      13'd1162: data <=16'b1111111110101100; 
      13'd1163: data <=16'b1111111101100011; 
      13'd1164: data <=16'b1111111111110111; 
      13'd1165: data <=16'b0000000010100111; 
      13'd1166: data <=16'b1111111110100001; 
      13'd1167: data <=16'b1111111111011110; 
      13'd1168: data <=16'b0000000000110010; 
      13'd1169: data <=16'b1111111110101001; 
      13'd1170: data <=16'b0000000011001010; 
      13'd1171: data <=16'b0000000000000110; 
      13'd1172: data <=16'b0000000000111011; 
      13'd1173: data <=16'b1111111110011101; 
      13'd1174: data <=16'b0000000000010011; 
      13'd1175: data <=16'b0000000010111100; 
      13'd1176: data <=16'b1111111111101110; 
      13'd1177: data <=16'b1111111110100000; 
      13'd1178: data <=16'b1111111110000001; 
      13'd1179: data <=16'b0000000000001000; 
      13'd1180: data <=16'b0000000000110010; 
      13'd1181: data <=16'b0000000001001110; 
      13'd1182: data <=16'b1111111110101000; 
      13'd1183: data <=16'b0000000000100011; 
      13'd1184: data <=16'b0000000010110011; 
      13'd1185: data <=16'b0000000001100101; 
      13'd1186: data <=16'b1111111110100111; 
      13'd1187: data <=16'b0000000001010101; 
      13'd1188: data <=16'b0000000000011111; 
      13'd1189: data <=16'b1111111110100000; 
      13'd1190: data <=16'b0000000001011000; 
      13'd1191: data <=16'b1111111101011011; 
      13'd1192: data <=16'b1111111110111101; 
      13'd1193: data <=16'b0000000010100111; 
      13'd1194: data <=16'b0000000000010001; 
      13'd1195: data <=16'b1111111110111100; 
      13'd1196: data <=16'b1111111110000100; 
      13'd1197: data <=16'b1111111111111010; 
      13'd1198: data <=16'b0000000011000010; 
      13'd1199: data <=16'b0000000000000011; 
      13'd1200: data <=16'b0000000001110010; 
      13'd1201: data <=16'b1111111111011111; 
      13'd1202: data <=16'b1111111101000011; 
      13'd1203: data <=16'b1111111111001101; 
      13'd1204: data <=16'b0000000010010011; 
      13'd1205: data <=16'b0000000010101111; 
      13'd1206: data <=16'b0000000001101110; 
      13'd1207: data <=16'b0000000000100000; 
      13'd1208: data <=16'b1111111111111001; 
      13'd1209: data <=16'b1111111111001110; 
      13'd1210: data <=16'b1111111110011010; 
      13'd1211: data <=16'b1111111110001001; 
      13'd1212: data <=16'b0000000001110001; 
      13'd1213: data <=16'b1111111111111010; 
      13'd1214: data <=16'b0000000001110100; 
      13'd1215: data <=16'b1111111110110110; 
      13'd1216: data <=16'b1111111110111100; 
      13'd1217: data <=16'b1111111111110101; 
      13'd1218: data <=16'b1111111111100111; 
      13'd1219: data <=16'b0000000000111100; 
      13'd1220: data <=16'b1111111110110000; 
      13'd1221: data <=16'b1111111111010110; 
      13'd1222: data <=16'b0000000001100001; 
      13'd1223: data <=16'b0000000001011100; 
      13'd1224: data <=16'b1111111110000000; 
      13'd1225: data <=16'b0000000001110101; 
      13'd1226: data <=16'b0000000000010001; 
      13'd1227: data <=16'b1111111111010100; 
      13'd1228: data <=16'b0000000000101110; 
      13'd1229: data <=16'b1111111100100000; 
      13'd1230: data <=16'b0000000000000011; 
      13'd1231: data <=16'b1111111111011110; 
      13'd1232: data <=16'b1111111111101000; 
      13'd1233: data <=16'b0000000001111001; 
      13'd1234: data <=16'b0000000000101011; 
      13'd1235: data <=16'b1111111110000001; 
      13'd1236: data <=16'b0000000000011000; 
      13'd1237: data <=16'b1111111111010100; 
      13'd1238: data <=16'b1111111110111101; 
      13'd1239: data <=16'b1111111110101001; 
      13'd1240: data <=16'b1111111111100110; 
      13'd1241: data <=16'b0000000000100100; 
      13'd1242: data <=16'b0000000000111101; 
      13'd1243: data <=16'b1111111101111000; 
      13'd1244: data <=16'b0000000000010101; 
      13'd1245: data <=16'b0000000001001111; 
      13'd1246: data <=16'b0000000001000101; 
      13'd1247: data <=16'b0000000000000111; 
      13'd1248: data <=16'b0000000001001010; 
      13'd1249: data <=16'b0000000010110000; 
      13'd1250: data <=16'b0000000001111010; 
      13'd1251: data <=16'b0000000000000110; 
      13'd1252: data <=16'b1111111111010101; 
      13'd1253: data <=16'b1111111111111100; 
      13'd1254: data <=16'b1111111111001011; 
      13'd1255: data <=16'b1111111111011100; 
      13'd1256: data <=16'b0000000001111001; 
      13'd1257: data <=16'b0000000001101010; 
      13'd1258: data <=16'b0000000001011100; 
      13'd1259: data <=16'b1111111100110001; 
      13'd1260: data <=16'b1111111111001000; 
      13'd1261: data <=16'b1111111110111010; 
      13'd1262: data <=16'b1111111111011001; 
      13'd1263: data <=16'b1111111111010000; 
      13'd1264: data <=16'b1111111111101110; 
      13'd1265: data <=16'b0000000010011011; 
      13'd1266: data <=16'b0000000000010011; 
      13'd1267: data <=16'b1111111110001011; 
      13'd1268: data <=16'b1111111101100111; 
      13'd1269: data <=16'b1111111111101011; 
      13'd1270: data <=16'b0000000001011101; 
      13'd1271: data <=16'b1111111111001111; 
      13'd1272: data <=16'b0000000000000110; 
      13'd1273: data <=16'b0000000000001010; 
      13'd1274: data <=16'b0000000000110000; 
      13'd1275: data <=16'b1111111111111001; 
      13'd1276: data <=16'b1111111111110011; 
      13'd1277: data <=16'b1111111110100111; 
      13'd1278: data <=16'b1111111111100111; 
      13'd1279: data <=16'b1111111111001000; 
      13'd1280: data <=16'b0000000000111011; 
      13'd1281: data <=16'b1111111111001011; 
      13'd1282: data <=16'b1111111110011111; 
      13'd1283: data <=16'b1111111110001100; 
      13'd1284: data <=16'b1111111110001011; 
      13'd1285: data <=16'b1111111111000000; 
      13'd1286: data <=16'b1111111111010001; 
      13'd1287: data <=16'b1111111111011110; 
      13'd1288: data <=16'b1111111111001110; 
      13'd1289: data <=16'b1111111101111111; 
      13'd1290: data <=16'b0000000000010001; 
      13'd1291: data <=16'b1111111101101111; 
      13'd1292: data <=16'b0000000001001000; 
      13'd1293: data <=16'b1111111111010000; 
      13'd1294: data <=16'b0000000001111000; 
      13'd1295: data <=16'b0000000001100110; 
      13'd1296: data <=16'b0000000010010100; 
      13'd1297: data <=16'b1111111110101110; 
      13'd1298: data <=16'b1111111111110001; 
      13'd1299: data <=16'b0000000000010011; 
      13'd1300: data <=16'b0000000000010110; 
      13'd1301: data <=16'b0000000000000000; 
      13'd1302: data <=16'b0000000000101111; 
      13'd1303: data <=16'b0000000010001010; 
      13'd1304: data <=16'b1111111111100010; 
      13'd1305: data <=16'b1111111111000001; 
      13'd1306: data <=16'b1111111110101010; 
      13'd1307: data <=16'b0000000000101100; 
      13'd1308: data <=16'b1111111111111010; 
      13'd1309: data <=16'b0000000001001101; 
      13'd1310: data <=16'b1111111110101010; 
      13'd1311: data <=16'b0000000010101100; 
      13'd1312: data <=16'b0000000010001111; 
      13'd1313: data <=16'b1111111111010110; 
      13'd1314: data <=16'b1111111110111001; 
      13'd1315: data <=16'b0000000000111100; 
      13'd1316: data <=16'b0000000000110111; 
      13'd1317: data <=16'b0000000000111001; 
      13'd1318: data <=16'b1111111110110010; 
      13'd1319: data <=16'b1111111100101011; 
      13'd1320: data <=16'b1111111111000010; 
      13'd1321: data <=16'b1111111101011011; 
      13'd1322: data <=16'b1111111110101100; 
      13'd1323: data <=16'b1111111110011010; 
      13'd1324: data <=16'b1111111110001100; 
      13'd1325: data <=16'b0000000000100100; 
      13'd1326: data <=16'b1111111101100001; 
      13'd1327: data <=16'b0000000001000110; 
      13'd1328: data <=16'b0000000001000111; 
      13'd1329: data <=16'b1111111111100100; 
      13'd1330: data <=16'b1111111101111001; 
      13'd1331: data <=16'b1111111111010011; 
      13'd1332: data <=16'b0000000000111001; 
      13'd1333: data <=16'b0000000000000001; 
      13'd1334: data <=16'b1111111100010001; 
      13'd1335: data <=16'b1111111111000101; 
      13'd1336: data <=16'b0000000010001010; 
      13'd1337: data <=16'b1111111111110000; 
      13'd1338: data <=16'b0000000010011000; 
      13'd1339: data <=16'b0000000000101111; 
      13'd1340: data <=16'b0000000001010011; 
      13'd1341: data <=16'b1111111111111101; 
      13'd1342: data <=16'b1111111111100101; 
      13'd1343: data <=16'b1111111111001110; 
      13'd1344: data <=16'b0000000010011010; 
      13'd1345: data <=16'b1111111111110000; 
      13'd1346: data <=16'b0000000001000111; 
      13'd1347: data <=16'b0000000000010011; 
      13'd1348: data <=16'b1111111111100000; 
      13'd1349: data <=16'b1111111101111011; 
      13'd1350: data <=16'b1111111111111111; 
      13'd1351: data <=16'b1111111111011001; 
      13'd1352: data <=16'b0000000000111011; 
      13'd1353: data <=16'b0000000000111110; 
      13'd1354: data <=16'b0000000010101011; 
      13'd1355: data <=16'b1111111111110100; 
      13'd1356: data <=16'b1111111110000000; 
      13'd1357: data <=16'b1111111111100100; 
      13'd1358: data <=16'b0000000000110001; 
      13'd1359: data <=16'b0000000000100001; 
      13'd1360: data <=16'b0000000000110111; 
      13'd1361: data <=16'b0000000000101100; 
      13'd1362: data <=16'b1111111111010111; 
      13'd1363: data <=16'b1111111100110100; 
      13'd1364: data <=16'b1111111111101100; 
      13'd1365: data <=16'b0000000000010010; 
      13'd1366: data <=16'b0000000011001110; 
      13'd1367: data <=16'b0000000001001010; 
      13'd1368: data <=16'b1111111111010011; 
      13'd1369: data <=16'b0000000000100110; 
      13'd1370: data <=16'b0000000000000001; 
      13'd1371: data <=16'b1111111111100110; 
      13'd1372: data <=16'b0000000000000000; 
      13'd1373: data <=16'b0000000001011001; 
      13'd1374: data <=16'b0000000000110100; 
      13'd1375: data <=16'b0000000000011111; 
      13'd1376: data <=16'b0000000011111111; 
      13'd1377: data <=16'b1111111110100000; 
      13'd1378: data <=16'b1111111110101001; 
      13'd1379: data <=16'b0000000010000101; 
      13'd1380: data <=16'b0000000000100111; 
      13'd1381: data <=16'b1111111111011111; 
      13'd1382: data <=16'b1111111111001000; 
      13'd1383: data <=16'b1111111110100111; 
      13'd1384: data <=16'b0000000000010010; 
      13'd1385: data <=16'b1111111111110100; 
      13'd1386: data <=16'b0000000000001010; 
      13'd1387: data <=16'b0000000000000000; 
      13'd1388: data <=16'b1111111111101101; 
      13'd1389: data <=16'b0000000000001101; 
      13'd1390: data <=16'b1111111110010110; 
      13'd1391: data <=16'b0000000010000110; 
      13'd1392: data <=16'b0000000010110101; 
      13'd1393: data <=16'b1111111111010101; 
      13'd1394: data <=16'b0000000000001010; 
      13'd1395: data <=16'b0000000000101100; 
      13'd1396: data <=16'b0000000000010001; 
      13'd1397: data <=16'b0000000010011111; 
      13'd1398: data <=16'b1111111110101110; 
      13'd1399: data <=16'b0000000010100001; 
      13'd1400: data <=16'b1111111110000001; 
      13'd1401: data <=16'b1111111110101101; 
      13'd1402: data <=16'b0000000000010011; 
      13'd1403: data <=16'b0000000000010011; 
      13'd1404: data <=16'b1111111110001011; 
      13'd1405: data <=16'b1111111101101001; 
      13'd1406: data <=16'b1111111111100001; 
      13'd1407: data <=16'b1111111110010001; 
      13'd1408: data <=16'b1111111101110001; 
      13'd1409: data <=16'b1111111111101100; 
      13'd1410: data <=16'b1111111110100110; 
      13'd1411: data <=16'b0000000000010110; 
      13'd1412: data <=16'b0000000000011111; 
      13'd1413: data <=16'b1111111110001001; 
      13'd1414: data <=16'b0000000000101010; 
      13'd1415: data <=16'b1111111101110001; 
      13'd1416: data <=16'b1111111101000001; 
      13'd1417: data <=16'b0000000000100001; 
      13'd1418: data <=16'b1111111110111011; 
      13'd1419: data <=16'b1111111100011111; 
      13'd1420: data <=16'b0000000010001101; 
      13'd1421: data <=16'b0000000000011100; 
      13'd1422: data <=16'b1111111111100000; 
      13'd1423: data <=16'b0000000000111110; 
      13'd1424: data <=16'b0000000000100011; 
      13'd1425: data <=16'b0000000001001100; 
      13'd1426: data <=16'b0000000001010111; 
      13'd1427: data <=16'b0000000000111011; 
      13'd1428: data <=16'b1111111111101010; 
      13'd1429: data <=16'b1111111111110111; 
      13'd1430: data <=16'b1111111111110110; 
      13'd1431: data <=16'b0000000010010011; 
      13'd1432: data <=16'b0000000000011011; 
      13'd1433: data <=16'b1111111111001010; 
      13'd1434: data <=16'b1111111110011011; 
      13'd1435: data <=16'b1111111101111100; 
      13'd1436: data <=16'b0000000000010001; 
      13'd1437: data <=16'b0000000001011010; 
      13'd1438: data <=16'b1111111111000100; 
      13'd1439: data <=16'b0000000000101010; 
      13'd1440: data <=16'b0000000001011100; 
      13'd1441: data <=16'b1111111101010001; 
      13'd1442: data <=16'b1111111111011000; 
      13'd1443: data <=16'b0000000000111101; 
      13'd1444: data <=16'b1111111111100011; 
      13'd1445: data <=16'b0000000001001000; 
      13'd1446: data <=16'b0000000010001011; 
      13'd1447: data <=16'b1111111111110111; 
      13'd1448: data <=16'b0000000000001000; 
      13'd1449: data <=16'b1111111111010010; 
      13'd1450: data <=16'b0000000010100000; 
      13'd1451: data <=16'b0000000000100010; 
      13'd1452: data <=16'b1111111110110110; 
      13'd1453: data <=16'b1111111110111000; 
      13'd1454: data <=16'b1111111110110111; 
      13'd1455: data <=16'b0000000011010011; 
      13'd1456: data <=16'b1111111110101101; 
      13'd1457: data <=16'b1111111110100010; 
      13'd1458: data <=16'b1111111111010111; 
      13'd1459: data <=16'b1111111110010111; 
      13'd1460: data <=16'b1111111111100011; 
      13'd1461: data <=16'b0000000001110100; 
      13'd1462: data <=16'b0000000001011101; 
      13'd1463: data <=16'b0000000001001101; 
      13'd1464: data <=16'b1111111111011111; 
      13'd1465: data <=16'b1111111111110011; 
      13'd1466: data <=16'b1111111110110010; 
      13'd1467: data <=16'b0000000001101000; 
      13'd1468: data <=16'b0000000000000010; 
      13'd1469: data <=16'b0000000000010110; 
      13'd1470: data <=16'b0000000000100100; 
      13'd1471: data <=16'b1111111110001100; 
      13'd1472: data <=16'b1111111100000010; 
      13'd1473: data <=16'b0000000001110001; 
      13'd1474: data <=16'b0000000001001110; 
      13'd1475: data <=16'b0000000000000110; 
      13'd1476: data <=16'b0000000010000110; 
      13'd1477: data <=16'b1111111111100010; 
      13'd1478: data <=16'b0000000010100111; 
      13'd1479: data <=16'b0000000010101011; 
      13'd1480: data <=16'b0000000000011111; 
      13'd1481: data <=16'b1111111111110111; 
      13'd1482: data <=16'b0000000010100110; 
      13'd1483: data <=16'b1111111110001010; 
      13'd1484: data <=16'b0000000000010100; 
      13'd1485: data <=16'b1111111110110010; 
      13'd1486: data <=16'b1111111111010110; 
      13'd1487: data <=16'b0000000001010101; 
      13'd1488: data <=16'b0000000000110001; 
      13'd1489: data <=16'b0000000000010001; 
      13'd1490: data <=16'b0000000001110010; 
      13'd1491: data <=16'b0000000000000101; 
      13'd1492: data <=16'b0000000000101100; 
      13'd1493: data <=16'b0000000000111100; 
      13'd1494: data <=16'b1111111111000001; 
      13'd1495: data <=16'b0000000001001101; 
      13'd1496: data <=16'b0000000000011100; 
      13'd1497: data <=16'b0000000000111111; 
      13'd1498: data <=16'b0000000001000011; 
      13'd1499: data <=16'b1111111110110000; 
      13'd1500: data <=16'b1111111111010001; 
      13'd1501: data <=16'b0000000100100011; 
      13'd1502: data <=16'b1111111110100110; 
      13'd1503: data <=16'b1111111111101001; 
      13'd1504: data <=16'b0000000001110110; 
      13'd1505: data <=16'b0000000001000010; 
      13'd1506: data <=16'b0000000000000010; 
      13'd1507: data <=16'b0000000001111110; 
      13'd1508: data <=16'b0000000000001001; 
      13'd1509: data <=16'b1111111111010011; 
      13'd1510: data <=16'b1111111110111110; 
      13'd1511: data <=16'b1111111111100111; 
      13'd1512: data <=16'b1111111111111000; 
      13'd1513: data <=16'b1111111111011110; 
      13'd1514: data <=16'b1111111110100100; 
      13'd1515: data <=16'b1111111110100111; 
      13'd1516: data <=16'b0000000010110011; 
      13'd1517: data <=16'b1111111111111010; 
      13'd1518: data <=16'b0000000000101010; 
      13'd1519: data <=16'b0000000000011010; 
      13'd1520: data <=16'b0000000010010010; 
      13'd1521: data <=16'b1111111110011010; 
      13'd1522: data <=16'b0000000000100001; 
      13'd1523: data <=16'b1111111101101011; 
      13'd1524: data <=16'b1111111111110011; 
      13'd1525: data <=16'b0000000001001101; 
      13'd1526: data <=16'b0000000001110010; 
      13'd1527: data <=16'b0000000000010011; 
      13'd1528: data <=16'b1111111111101100; 
      13'd1529: data <=16'b0000000001011011; 
      13'd1530: data <=16'b0000000000101000; 
      13'd1531: data <=16'b1111111101000001; 
      13'd1532: data <=16'b1111111110110001; 
      13'd1533: data <=16'b1111111111010010; 
      13'd1534: data <=16'b0000000001100001; 
      13'd1535: data <=16'b0000000001110101; 
      13'd1536: data <=16'b0000000001010001; 
      13'd1537: data <=16'b1111111110101000; 
      13'd1538: data <=16'b0000000001001010; 
      13'd1539: data <=16'b1111111111111111; 
      13'd1540: data <=16'b0000000010001101; 
      13'd1541: data <=16'b1111111111101111; 
      13'd1542: data <=16'b0000000010101011; 
      13'd1543: data <=16'b1111111101111110; 
      13'd1544: data <=16'b1111111111110100; 
      13'd1545: data <=16'b1111111111110010; 
      13'd1546: data <=16'b1111111110100111; 
      13'd1547: data <=16'b0000000000100011; 
      13'd1548: data <=16'b1111111111000101; 
      13'd1549: data <=16'b1111111111100010; 
      13'd1550: data <=16'b0000000001011110; 
      13'd1551: data <=16'b0000000001011111; 
      13'd1552: data <=16'b0000000000001111; 
      13'd1553: data <=16'b1111111111010000; 
      13'd1554: data <=16'b1111111111000100; 
      13'd1555: data <=16'b1111111111001001; 
      13'd1556: data <=16'b0000000000110011; 
      13'd1557: data <=16'b0000000001101010; 
      13'd1558: data <=16'b1111111111111000; 
      13'd1559: data <=16'b0000000000100101; 
      13'd1560: data <=16'b0000000000110000; 
      13'd1561: data <=16'b0000000000001010; 
      13'd1562: data <=16'b0000000000101111; 
      13'd1563: data <=16'b0000000010001101; 
      13'd1564: data <=16'b1111111101001100; 
      13'd1565: data <=16'b0000000001010101; 
      13'd1566: data <=16'b1111111101110000; 
      13'd1567: data <=16'b1111111101001000; 
      13'd1568: data <=16'b1111111101011011; 
      13'd1569: data <=16'b0000000001110011; 
      13'd1570: data <=16'b0000000001110101; 
      13'd1571: data <=16'b1111111110001011; 
      13'd1572: data <=16'b0000000000011101; 
      13'd1573: data <=16'b1111111111000110; 
      13'd1574: data <=16'b0000000000001100; 
      13'd1575: data <=16'b1111111110110100; 
      13'd1576: data <=16'b1111111110111100; 
      13'd1577: data <=16'b1111111111011000; 
      13'd1578: data <=16'b1111111110100011; 
      13'd1579: data <=16'b1111111110010100; 
      13'd1580: data <=16'b0000000000101011; 
      13'd1581: data <=16'b0000000000100110; 
      13'd1582: data <=16'b0000000000001100; 
      13'd1583: data <=16'b0000000000001111; 
      13'd1584: data <=16'b0000000000111000; 
      13'd1585: data <=16'b1111111111010111; 
      13'd1586: data <=16'b0000000001100100; 
      13'd1587: data <=16'b0000000000010001; 
      13'd1588: data <=16'b0000000000001000; 
      13'd1589: data <=16'b0000000000110111; 
      13'd1590: data <=16'b0000000001100110; 
      13'd1591: data <=16'b1111111111000010; 
      13'd1592: data <=16'b1111111110000011; 
      13'd1593: data <=16'b1111111111111010; 
      13'd1594: data <=16'b0000000001111001; 
      13'd1595: data <=16'b0000000000101010; 
      13'd1596: data <=16'b0000000100000011; 
      13'd1597: data <=16'b1111111110010001; 
      13'd1598: data <=16'b1111111110010010; 
      13'd1599: data <=16'b1111111110101100; 
      13'd1600: data <=16'b1111111111000011; 
      13'd1601: data <=16'b1111111101001100; 
      13'd1602: data <=16'b0000000000101001; 
      13'd1603: data <=16'b0000000000110000; 
      13'd1604: data <=16'b0000000010100001; 
      13'd1605: data <=16'b1111111110001010; 
      13'd1606: data <=16'b1111111111000000; 
      13'd1607: data <=16'b0000000000100101; 
      13'd1608: data <=16'b1111111110100101; 
      13'd1609: data <=16'b0000000000011001; 
      13'd1610: data <=16'b0000000010001010; 
      13'd1611: data <=16'b0000000001010011; 
      13'd1612: data <=16'b1111111110001100; 
      13'd1613: data <=16'b0000000000011110; 
      13'd1614: data <=16'b0000000001010010; 
      13'd1615: data <=16'b0000000001101000; 
      13'd1616: data <=16'b0000000000101110; 
      13'd1617: data <=16'b0000000010110100; 
      13'd1618: data <=16'b0000000001000000; 
      13'd1619: data <=16'b0000000000111000; 
      13'd1620: data <=16'b1111111110110011; 
      13'd1621: data <=16'b0000000000110101; 
      13'd1622: data <=16'b0000000011000010; 
      13'd1623: data <=16'b0000000001110000; 
      13'd1624: data <=16'b1111111110110111; 
      13'd1625: data <=16'b0000000000010110; 
      13'd1626: data <=16'b0000000000010000; 
      13'd1627: data <=16'b0000000000011010; 
      13'd1628: data <=16'b1111111111010001; 
      13'd1629: data <=16'b0000000000101100; 
      13'd1630: data <=16'b1111111110110000; 
      13'd1631: data <=16'b1111111111010010; 
      13'd1632: data <=16'b0000000010001010; 
      13'd1633: data <=16'b1111111111011010; 
      13'd1634: data <=16'b1111111110101110; 
      13'd1635: data <=16'b0000000010110011; 
      13'd1636: data <=16'b0000000010000100; 
      13'd1637: data <=16'b1111111111000111; 
      13'd1638: data <=16'b0000000001000011; 
      13'd1639: data <=16'b0000000000001011; 
      13'd1640: data <=16'b1111111100000001; 
      13'd1641: data <=16'b0000000001000001; 
      13'd1642: data <=16'b1111111110111000; 
      13'd1643: data <=16'b1111111111101011; 
      13'd1644: data <=16'b0000000001100101; 
      13'd1645: data <=16'b0000000000011111; 
      13'd1646: data <=16'b0000000000100000; 
      13'd1647: data <=16'b0000000001110110; 
      13'd1648: data <=16'b1111111111110101; 
      13'd1649: data <=16'b1111111111000111; 
      13'd1650: data <=16'b1111111111000000; 
      13'd1651: data <=16'b0000000000001010; 
      13'd1652: data <=16'b1111111111010011; 
      13'd1653: data <=16'b0000000001010000; 
      13'd1654: data <=16'b1111111110100111; 
      13'd1655: data <=16'b1111111110000011; 
      13'd1656: data <=16'b0000000000000011; 
      13'd1657: data <=16'b1111111110000111; 
      13'd1658: data <=16'b1111111110000110; 
      13'd1659: data <=16'b1111111110111111; 
      13'd1660: data <=16'b1111111110111100; 
      13'd1661: data <=16'b0000000000100111; 
      13'd1662: data <=16'b1111111111110011; 
      13'd1663: data <=16'b1111111110100000; 
      13'd1664: data <=16'b0000000000111110; 
      13'd1665: data <=16'b0000000000111011; 
      13'd1666: data <=16'b1111111110101010; 
      13'd1667: data <=16'b1111111111100000; 
      13'd1668: data <=16'b1111111110000100; 
      13'd1669: data <=16'b1111111110101111; 
      13'd1670: data <=16'b1111111110100010; 
      13'd1671: data <=16'b0000000001111010; 
      13'd1672: data <=16'b1111111111101010; 
      13'd1673: data <=16'b1111111111111001; 
      13'd1674: data <=16'b1111111110011110; 
      13'd1675: data <=16'b0000000001000101; 
      13'd1676: data <=16'b0000000001011011; 
      13'd1677: data <=16'b0000000000100101; 
      13'd1678: data <=16'b1111111110000010; 
      13'd1679: data <=16'b0000000000001100; 
      13'd1680: data <=16'b1111111100101100; 
      13'd1681: data <=16'b1111111111100101; 
      13'd1682: data <=16'b0000000000110000; 
      13'd1683: data <=16'b0000000000001101; 
      13'd1684: data <=16'b1111111111101110; 
      13'd1685: data <=16'b0000000000111110; 
      13'd1686: data <=16'b1111111110000010; 
      13'd1687: data <=16'b0000000000011111; 
      13'd1688: data <=16'b1111111111111011; 
      13'd1689: data <=16'b0000000000011110; 
      13'd1690: data <=16'b0000000000110100; 
      13'd1691: data <=16'b0000000001000110; 
      13'd1692: data <=16'b0000000000010011; 
      13'd1693: data <=16'b1111111110010000; 
      13'd1694: data <=16'b1111111111011010; 
      13'd1695: data <=16'b1111111111011111; 
      13'd1696: data <=16'b1111111111110111; 
      13'd1697: data <=16'b0000000001000001; 
      13'd1698: data <=16'b0000000001001011; 
      13'd1699: data <=16'b0000000000010100; 
      13'd1700: data <=16'b1111111110011111; 
      13'd1701: data <=16'b1111111110100110; 
      13'd1702: data <=16'b0000000011101110; 
      13'd1703: data <=16'b1111111101101111; 
      13'd1704: data <=16'b0000000000010111; 
      13'd1705: data <=16'b0000000000101100; 
      13'd1706: data <=16'b0000000010000000; 
      13'd1707: data <=16'b0000000000010101; 
      13'd1708: data <=16'b1111111110110010; 
      13'd1709: data <=16'b0000000001000011; 
      13'd1710: data <=16'b0000000000111001; 
      13'd1711: data <=16'b1111111111111101; 
      13'd1712: data <=16'b0000000000011111; 
      13'd1713: data <=16'b1111111110111101; 
      13'd1714: data <=16'b1111111110010001; 
      13'd1715: data <=16'b1111111111010111; 
      13'd1716: data <=16'b0000000011010000; 
      13'd1717: data <=16'b0000000001101110; 
      13'd1718: data <=16'b0000000000010010; 
      13'd1719: data <=16'b1111111111101110; 
      13'd1720: data <=16'b1111111111011001; 
      13'd1721: data <=16'b0000000000011100; 
      13'd1722: data <=16'b0000000001010000; 
      13'd1723: data <=16'b0000000001011101; 
      13'd1724: data <=16'b0000000000010010; 
      13'd1725: data <=16'b1111111101101101; 
      13'd1726: data <=16'b0000000000100010; 
      13'd1727: data <=16'b0000000000011010; 
      13'd1728: data <=16'b1111111101101110; 
      13'd1729: data <=16'b0000000010011110; 
      13'd1730: data <=16'b0000000010000000; 
      13'd1731: data <=16'b1111111110010011; 
      13'd1732: data <=16'b0000000000010100; 
      13'd1733: data <=16'b1111111110011101; 
      13'd1734: data <=16'b0000000000101011; 
      13'd1735: data <=16'b0000000000011100; 
      13'd1736: data <=16'b0000000000011010; 
      13'd1737: data <=16'b1111111111111010; 
      13'd1738: data <=16'b0000000000001110; 
      13'd1739: data <=16'b1111111110100000; 
      13'd1740: data <=16'b0000000001001111; 
      13'd1741: data <=16'b0000000001101001; 
      13'd1742: data <=16'b0000000001000101; 
      13'd1743: data <=16'b1111111110101100; 
      13'd1744: data <=16'b1111111110001010; 
      13'd1745: data <=16'b1111111111101111; 
      13'd1746: data <=16'b1111111110101010; 
      13'd1747: data <=16'b0000000000111101; 
      13'd1748: data <=16'b1111111111110001; 
      13'd1749: data <=16'b0000000011100101; 
      13'd1750: data <=16'b0000000000001011; 
      13'd1751: data <=16'b0000000000100001; 
      13'd1752: data <=16'b0000000010001011; 
      13'd1753: data <=16'b1111111111001010; 
      13'd1754: data <=16'b1111111110011101; 
      13'd1755: data <=16'b1111111111110000; 
      13'd1756: data <=16'b0000000000000000; 
      13'd1757: data <=16'b1111111110110000; 
      13'd1758: data <=16'b1111111111000011; 
      13'd1759: data <=16'b0000000001101000; 
      13'd1760: data <=16'b0000000000010100; 
      13'd1761: data <=16'b0000000001000000; 
      13'd1762: data <=16'b1111111110111011; 
      13'd1763: data <=16'b0000000000001001; 
      13'd1764: data <=16'b0000000000111101; 
      13'd1765: data <=16'b1111111110001111; 
      13'd1766: data <=16'b1111111111100101; 
      13'd1767: data <=16'b0000000010000101; 
      13'd1768: data <=16'b1111111111000001; 
      13'd1769: data <=16'b0000000000110000; 
      13'd1770: data <=16'b1111111111111100; 
      13'd1771: data <=16'b1111111011010101; 
      13'd1772: data <=16'b0000000001011010; 
      13'd1773: data <=16'b1111111101010011; 
      13'd1774: data <=16'b0000000000111100; 
      13'd1775: data <=16'b0000000010110011; 
      13'd1776: data <=16'b1111111110101011; 
      13'd1777: data <=16'b1111111111000001; 
      13'd1778: data <=16'b0000000010000100; 
      13'd1779: data <=16'b1111111111100101; 
      13'd1780: data <=16'b1111111111110001; 
      13'd1781: data <=16'b0000000010011011; 
      13'd1782: data <=16'b0000000010001000; 
      13'd1783: data <=16'b0000000000101101; 
      13'd1784: data <=16'b1111111101010100; 
      13'd1785: data <=16'b1111111110010011; 
      13'd1786: data <=16'b1111111110011000; 
      13'd1787: data <=16'b1111111101011110; 
      13'd1788: data <=16'b0000000000001110; 
      13'd1789: data <=16'b0000000001111101; 
      13'd1790: data <=16'b1111111101100110; 
      13'd1791: data <=16'b0000000000110000; 
      13'd1792: data <=16'b0000000000011111; 
      13'd1793: data <=16'b1111111111001100; 
      13'd1794: data <=16'b1111111110111100; 
      13'd1795: data <=16'b1111111111111101; 
      13'd1796: data <=16'b0000000001111100; 
      13'd1797: data <=16'b1111111111111010; 
      13'd1798: data <=16'b0000000010010011; 
      13'd1799: data <=16'b0000000000100100; 
      13'd1800: data <=16'b1111111111101001; 
      13'd1801: data <=16'b1111111101000010; 
      13'd1802: data <=16'b0000000000001001; 
      13'd1803: data <=16'b1111111111000011; 
      13'd1804: data <=16'b0000000000110110; 
      13'd1805: data <=16'b0000000010000101; 
      13'd1806: data <=16'b0000000000011010; 
      13'd1807: data <=16'b0000000010010010; 
      13'd1808: data <=16'b1111111101110110; 
      13'd1809: data <=16'b1111111110100110; 
      13'd1810: data <=16'b0000000000010111; 
      13'd1811: data <=16'b1111111111110111; 
      13'd1812: data <=16'b1111111111111101; 
      13'd1813: data <=16'b0000000000000101; 
      13'd1814: data <=16'b0000000000011111; 
      13'd1815: data <=16'b0000000000100011; 
      13'd1816: data <=16'b0000000010001001; 
      13'd1817: data <=16'b0000000001000010; 
      13'd1818: data <=16'b0000000010111011; 
      13'd1819: data <=16'b1111111111101010; 
      13'd1820: data <=16'b1111111101111001; 
      13'd1821: data <=16'b1111111111010111; 
      13'd1822: data <=16'b1111111110100010; 
      13'd1823: data <=16'b0000000000101001; 
      13'd1824: data <=16'b0000000000000111; 
      13'd1825: data <=16'b1111111101111111; 
      13'd1826: data <=16'b1111111110001100; 
      13'd1827: data <=16'b1111111111100011; 
      13'd1828: data <=16'b0000000000001011; 
      13'd1829: data <=16'b1111111111010001; 
      13'd1830: data <=16'b0000000001001010; 
      13'd1831: data <=16'b1111111111110110; 
      13'd1832: data <=16'b0000000000101111; 
      13'd1833: data <=16'b1111111111100110; 
      13'd1834: data <=16'b0000000000101110; 
      13'd1835: data <=16'b0000000001001110; 
      13'd1836: data <=16'b0000000001100101; 
      13'd1837: data <=16'b0000000000011001; 
      13'd1838: data <=16'b0000000000001011; 
      13'd1839: data <=16'b1111111110001111; 
      13'd1840: data <=16'b0000000010000110; 
      13'd1841: data <=16'b0000000001011010; 
      13'd1842: data <=16'b1111111111001010; 
      13'd1843: data <=16'b1111111110110111; 
      13'd1844: data <=16'b1111111110110111; 
      13'd1845: data <=16'b1111111111100101; 
      13'd1846: data <=16'b1111111100111111; 
      13'd1847: data <=16'b0000000000011001; 
      13'd1848: data <=16'b0000000000100111; 
      13'd1849: data <=16'b1111111111011100; 
      13'd1850: data <=16'b0000000001101000; 
      13'd1851: data <=16'b0000000010000100; 
      13'd1852: data <=16'b0000000001010100; 
      13'd1853: data <=16'b0000000000111000; 
      13'd1854: data <=16'b1111111101001000; 
      13'd1855: data <=16'b0000000000111011; 
      13'd1856: data <=16'b1111111111010011; 
      13'd1857: data <=16'b1111111111010101; 
      13'd1858: data <=16'b0000000010010010; 
      13'd1859: data <=16'b0000000001110011; 
      13'd1860: data <=16'b1111111110110100; 
      13'd1861: data <=16'b1111111111010001; 
      13'd1862: data <=16'b0000000000000010; 
      13'd1863: data <=16'b0000000000111101; 
      13'd1864: data <=16'b0000000000101001; 
      13'd1865: data <=16'b0000000000101000; 
      13'd1866: data <=16'b1111111111101011; 
      13'd1867: data <=16'b0000000001010010; 
      13'd1868: data <=16'b1111111110011100; 
      13'd1869: data <=16'b0000000000110101; 
      13'd1870: data <=16'b1111111111010000; 
      13'd1871: data <=16'b1111111111100000; 
      13'd1872: data <=16'b1111111101001100; 
      13'd1873: data <=16'b0000000000000100; 
      13'd1874: data <=16'b0000000001010100; 
      13'd1875: data <=16'b1111111111100010; 
      13'd1876: data <=16'b1111111100001111; 
      13'd1877: data <=16'b0000000011001010; 
      13'd1878: data <=16'b0000000000110101; 
      13'd1879: data <=16'b1111111111101101; 
      13'd1880: data <=16'b0000000000010101; 
      13'd1881: data <=16'b0000000000001000; 
      13'd1882: data <=16'b0000000000010101; 
      13'd1883: data <=16'b0000000001001011; 
      13'd1884: data <=16'b0000000000111010; 
      13'd1885: data <=16'b1111111101110101; 
      13'd1886: data <=16'b1111111101110100; 
      13'd1887: data <=16'b1111111101011001; 
      13'd1888: data <=16'b1111111111100011; 
      13'd1889: data <=16'b1111111101111010; 
      13'd1890: data <=16'b1111111111110010; 
      13'd1891: data <=16'b1111111110110100; 
      13'd1892: data <=16'b0000000000100011; 
      13'd1893: data <=16'b0000000000010110; 
      13'd1894: data <=16'b0000000010100100; 
      13'd1895: data <=16'b1111111111000110; 
      13'd1896: data <=16'b1111111110011111; 
      13'd1897: data <=16'b1111111100111101; 
      13'd1898: data <=16'b0000000000011001; 
      13'd1899: data <=16'b1111111111110110; 
      13'd1900: data <=16'b1111111110010101; 
      13'd1901: data <=16'b0000000000100100; 
      13'd1902: data <=16'b1111111111100001; 
      13'd1903: data <=16'b0000000000110010; 
      13'd1904: data <=16'b0000000000001001; 
      13'd1905: data <=16'b1111111110101000; 
      13'd1906: data <=16'b0000000010110000; 
      13'd1907: data <=16'b1111111101110101; 
      13'd1908: data <=16'b0000000001000011; 
      13'd1909: data <=16'b1111111111101011; 
      13'd1910: data <=16'b1111111101101110; 
      13'd1911: data <=16'b0000000010010010; 
      13'd1912: data <=16'b1111111111111011; 
      13'd1913: data <=16'b1111111111000101; 
      13'd1914: data <=16'b1111111110001001; 
      13'd1915: data <=16'b1111111111011110; 
      13'd1916: data <=16'b1111111110100000; 
      13'd1917: data <=16'b1111111110100110; 
      13'd1918: data <=16'b0000000001010111; 
      13'd1919: data <=16'b1111111111101011; 
      13'd1920: data <=16'b0000000010011100; 
      13'd1921: data <=16'b0000000010110011; 
      13'd1922: data <=16'b1111111111011001; 
      13'd1923: data <=16'b0000000000000011; 
      13'd1924: data <=16'b0000000001000101; 
      13'd1925: data <=16'b1111111111011100; 
      13'd1926: data <=16'b1111111110101110; 
      13'd1927: data <=16'b0000000001100001; 
      13'd1928: data <=16'b1111111101111101; 
      13'd1929: data <=16'b0000000000100010; 
      13'd1930: data <=16'b1111111110100100; 
      13'd1931: data <=16'b1111111110111000; 
      13'd1932: data <=16'b0000000000111000; 
      13'd1933: data <=16'b1111111011101010; 
      13'd1934: data <=16'b1111111110010101; 
      13'd1935: data <=16'b1111111111000101; 
      13'd1936: data <=16'b1111111110111110; 
      13'd1937: data <=16'b0000000000100111; 
      13'd1938: data <=16'b1111111110111100; 
      13'd1939: data <=16'b1111111111000001; 
      13'd1940: data <=16'b1111111111000110; 
      13'd1941: data <=16'b0000000000000111; 
      13'd1942: data <=16'b1111111110100010; 
      13'd1943: data <=16'b0000000000001110; 
      13'd1944: data <=16'b1111111111100011; 
      13'd1945: data <=16'b0000000001111111; 
      13'd1946: data <=16'b0000000001000011; 
      13'd1947: data <=16'b1111111110000011; 
      13'd1948: data <=16'b0000000010111100; 
      13'd1949: data <=16'b0000000000011010; 
      13'd1950: data <=16'b1111111101110100; 
      13'd1951: data <=16'b1111111111001010; 
      13'd1952: data <=16'b1111111110111110; 
      13'd1953: data <=16'b1111111110101000; 
      13'd1954: data <=16'b0000000000100000; 
      13'd1955: data <=16'b0000000010000011; 
      13'd1956: data <=16'b0000000010100100; 
      13'd1957: data <=16'b0000000000011000; 
      13'd1958: data <=16'b0000000011000001; 
      13'd1959: data <=16'b1111111110110101; 
      13'd1960: data <=16'b1111111101111000; 
      13'd1961: data <=16'b0000000001001000; 
      13'd1962: data <=16'b1111111111100110; 
      13'd1963: data <=16'b1111111111111100; 
      13'd1964: data <=16'b1111111110100110; 
      13'd1965: data <=16'b0000000001100001; 
      13'd1966: data <=16'b1111111111100110; 
      13'd1967: data <=16'b0000000001001011; 
      13'd1968: data <=16'b1111111111000100; 
      13'd1969: data <=16'b0000000010010100; 
      13'd1970: data <=16'b1111111111101001; 
      13'd1971: data <=16'b0000000001001100; 
      13'd1972: data <=16'b1111111110000100; 
      13'd1973: data <=16'b0000000011000010; 
      13'd1974: data <=16'b0000000000111111; 
      13'd1975: data <=16'b0000000001000101; 
      13'd1976: data <=16'b1111111110101101; 
      13'd1977: data <=16'b0000000000111101; 
      13'd1978: data <=16'b1111111111000000; 
      13'd1979: data <=16'b1111111110111100; 
      13'd1980: data <=16'b1111111110101010; 
      13'd1981: data <=16'b1111111101111111; 
      13'd1982: data <=16'b1111111111001010; 
      13'd1983: data <=16'b1111111110110111; 
      13'd1984: data <=16'b0000000000111100; 
      13'd1985: data <=16'b0000000000011000; 
      13'd1986: data <=16'b0000000000101000; 
      13'd1987: data <=16'b0000000001010000; 
      13'd1988: data <=16'b1111111111001100; 
      13'd1989: data <=16'b1111111111100011; 
      13'd1990: data <=16'b0000000010100111; 
      13'd1991: data <=16'b0000000000000110; 
      13'd1992: data <=16'b0000000000001011; 
      13'd1993: data <=16'b0000000000110101; 
      13'd1994: data <=16'b0000000001000011; 
      13'd1995: data <=16'b0000000001111000; 
      13'd1996: data <=16'b0000000000110101; 
      13'd1997: data <=16'b1111111111001010; 
      13'd1998: data <=16'b0000000001010010; 
      13'd1999: data <=16'b0000000000011111; 
      13'd2000: data <=16'b1111111111101101; 
      13'd2001: data <=16'b1111111111111111; 
      13'd2002: data <=16'b0000000000010111; 
      13'd2003: data <=16'b0000000001010111; 
      13'd2004: data <=16'b0000000000001000; 
      13'd2005: data <=16'b0000000000011000; 
      13'd2006: data <=16'b1111111110000000; 
      13'd2007: data <=16'b0000000000100011; 
      13'd2008: data <=16'b0000000000100010; 
      13'd2009: data <=16'b0000000010001000; 
      13'd2010: data <=16'b0000000000100110; 
      13'd2011: data <=16'b1111111110011110; 
      13'd2012: data <=16'b0000000001001000; 
      13'd2013: data <=16'b0000000000001111; 
      13'd2014: data <=16'b0000000001001101; 
      13'd2015: data <=16'b0000000001010100; 
      13'd2016: data <=16'b0000000011101110; 
      13'd2017: data <=16'b0000000001110010; 
      13'd2018: data <=16'b1111111101101011; 
      13'd2019: data <=16'b0000000000110000; 
      13'd2020: data <=16'b1111111111101111; 
      13'd2021: data <=16'b1111111110100000; 
      13'd2022: data <=16'b1111111110010100; 
      13'd2023: data <=16'b1111111111000011; 
      13'd2024: data <=16'b1111111111001100; 
      13'd2025: data <=16'b0000000000001101; 
      13'd2026: data <=16'b1111111111000110; 
      13'd2027: data <=16'b1111111111101111; 
      13'd2028: data <=16'b0000000000011110; 
      13'd2029: data <=16'b0000000000010110; 
      13'd2030: data <=16'b0000000000001110; 
      13'd2031: data <=16'b0000000010001011; 
      13'd2032: data <=16'b0000000001011111; 
      13'd2033: data <=16'b0000000000111111; 
      13'd2034: data <=16'b0000000000010010; 
      13'd2035: data <=16'b0000000001000010; 
      13'd2036: data <=16'b1111111111111001; 
      13'd2037: data <=16'b0000000001001001; 
      13'd2038: data <=16'b1111111111000110; 
      13'd2039: data <=16'b1111111111101110; 
      13'd2040: data <=16'b0000000001000100; 
      13'd2041: data <=16'b1111111101100101; 
      13'd2042: data <=16'b1111111111110100; 
      13'd2043: data <=16'b0000000001000111; 
      13'd2044: data <=16'b0000000000110000; 
      13'd2045: data <=16'b0000000011011111; 
      13'd2046: data <=16'b1111111110101010; 
      13'd2047: data <=16'b0000000001001001; 
      13'd2048: data <=16'b1111111111010010; 
      13'd2049: data <=16'b0000000000000010; 
      13'd2050: data <=16'b1111111110001011; 
      13'd2051: data <=16'b0000000000111010; 
      13'd2052: data <=16'b1111111111110000; 
      13'd2053: data <=16'b1111111111011000; 
      13'd2054: data <=16'b0000000001111101; 
      13'd2055: data <=16'b1111111100100111; 
      13'd2056: data <=16'b1111111111100000; 
      13'd2057: data <=16'b1111111110011001; 
      13'd2058: data <=16'b0000000000100110; 
      13'd2059: data <=16'b0000000010001000; 
      13'd2060: data <=16'b0000000000000110; 
      13'd2061: data <=16'b0000000000011001; 
      13'd2062: data <=16'b1111111110000000; 
      13'd2063: data <=16'b0000000001101000; 
      13'd2064: data <=16'b1111111111100010; 
      13'd2065: data <=16'b0000000000110010; 
      13'd2066: data <=16'b1111111110101001; 
      13'd2067: data <=16'b1111111111001001; 
      13'd2068: data <=16'b0000000001111111; 
      13'd2069: data <=16'b0000000000101011; 
      13'd2070: data <=16'b1111111100110001; 
      13'd2071: data <=16'b1111111111110000; 
      13'd2072: data <=16'b0000000000010111; 
      13'd2073: data <=16'b0000000001111011; 
      13'd2074: data <=16'b0000000001001111; 
      13'd2075: data <=16'b0000000010001100; 
      13'd2076: data <=16'b1111111101001100; 
      13'd2077: data <=16'b1111111111010001; 
      13'd2078: data <=16'b0000000001000000; 
      13'd2079: data <=16'b0000000001110111; 
      13'd2080: data <=16'b0000000000010101; 
      13'd2081: data <=16'b1111111110100010; 
      13'd2082: data <=16'b0000000011010001; 
      13'd2083: data <=16'b0000000000000010; 
      13'd2084: data <=16'b0000000000001000; 
      13'd2085: data <=16'b0000000010001011; 
      13'd2086: data <=16'b1111111110010101; 
      13'd2087: data <=16'b0000000000101111; 
      13'd2088: data <=16'b0000000001001000; 
      13'd2089: data <=16'b1111111101010000; 
      13'd2090: data <=16'b1111111110101101; 
      13'd2091: data <=16'b1111111111001101; 
      13'd2092: data <=16'b0000000001100011; 
      13'd2093: data <=16'b1111111111001100; 
      13'd2094: data <=16'b1111111111101110; 
      13'd2095: data <=16'b1111111100111010; 
      13'd2096: data <=16'b0000000001111011; 
      13'd2097: data <=16'b1111111111101010; 
      13'd2098: data <=16'b0000000000011000; 
      13'd2099: data <=16'b1111111110101001; 
      13'd2100: data <=16'b0000000001010011; 
      13'd2101: data <=16'b1111111110110110; 
      13'd2102: data <=16'b0000000001011100; 
      13'd2103: data <=16'b1111111111010110; 
      13'd2104: data <=16'b0000000000001000; 
      13'd2105: data <=16'b1111111111110000; 
      13'd2106: data <=16'b0000000000001111; 
      13'd2107: data <=16'b0000000010110110; 
      13'd2108: data <=16'b1111111111100111; 
      13'd2109: data <=16'b0000000000111001; 
      13'd2110: data <=16'b0000000000001000; 
      13'd2111: data <=16'b1111111111010001; 
      13'd2112: data <=16'b1111111101110011; 
      13'd2113: data <=16'b1111111110110110; 
      13'd2114: data <=16'b1111111110100001; 
      13'd2115: data <=16'b0000000000011100; 
      13'd2116: data <=16'b1111111110110110; 
      13'd2117: data <=16'b1111111110110100; 
      13'd2118: data <=16'b0000000001001001; 
      13'd2119: data <=16'b1111111111111100; 
      13'd2120: data <=16'b0000000000011010; 
      13'd2121: data <=16'b1111111111001101; 
      13'd2122: data <=16'b0000000000100001; 
      13'd2123: data <=16'b0000000000101011; 
      13'd2124: data <=16'b0000000001000000; 
      13'd2125: data <=16'b0000000010000000; 
      13'd2126: data <=16'b0000000001001110; 
      13'd2127: data <=16'b1111111111100011; 
      13'd2128: data <=16'b0000000001001111; 
      13'd2129: data <=16'b1111111110011100; 
      13'd2130: data <=16'b1111111110101111; 
      13'd2131: data <=16'b1111111111011001; 
      13'd2132: data <=16'b1111111101110011; 
      13'd2133: data <=16'b1111111111100101; 
      13'd2134: data <=16'b1111111110110000; 
      13'd2135: data <=16'b0000000001011110; 
      13'd2136: data <=16'b1111111101111000; 
      13'd2137: data <=16'b0000000000101011; 
      13'd2138: data <=16'b1111111111011111; 
      13'd2139: data <=16'b0000000000110111; 
      13'd2140: data <=16'b1111111111111100; 
      13'd2141: data <=16'b1111111111000000; 
      13'd2142: data <=16'b0000000001100011; 
      13'd2143: data <=16'b1111111101100101; 
      13'd2144: data <=16'b0000000010011011; 
      13'd2145: data <=16'b1111111101001101; 
      13'd2146: data <=16'b1111111111101110; 
      13'd2147: data <=16'b1111111100001100; 
      13'd2148: data <=16'b1111111110011010; 
      13'd2149: data <=16'b0000000010100010; 
      13'd2150: data <=16'b0000000000000010; 
      13'd2151: data <=16'b0000000010100011; 
      13'd2152: data <=16'b0000000000110010; 
      13'd2153: data <=16'b1111111101011001; 
      13'd2154: data <=16'b1111111111110111; 
      13'd2155: data <=16'b0000000000110100; 
      13'd2156: data <=16'b1111111101000110; 
      13'd2157: data <=16'b1111111111101000; 
      13'd2158: data <=16'b1111111111010101; 
      13'd2159: data <=16'b0000000001001011; 
      13'd2160: data <=16'b1111111110010100; 
      13'd2161: data <=16'b0000000001100101; 
      13'd2162: data <=16'b1111111111111001; 
      13'd2163: data <=16'b1111111101011111; 
      13'd2164: data <=16'b0000000000101010; 
      13'd2165: data <=16'b1111111101010101; 
      13'd2166: data <=16'b0000000000001010; 
      13'd2167: data <=16'b0000000000110000; 
      13'd2168: data <=16'b0000000000110011; 
      13'd2169: data <=16'b1111111101111101; 
      13'd2170: data <=16'b1111111111100100; 
      13'd2171: data <=16'b0000000000111001; 
      13'd2172: data <=16'b1111111110000110; 
      13'd2173: data <=16'b1111111111010110; 
      13'd2174: data <=16'b0000000001011011; 
      13'd2175: data <=16'b1111111111000101; 
      13'd2176: data <=16'b0000000000000010; 
      13'd2177: data <=16'b1111111111110111; 
      13'd2178: data <=16'b0000000010001101; 
      13'd2179: data <=16'b1111111100101010; 
      13'd2180: data <=16'b1111111110111111; 
      13'd2181: data <=16'b1111111111010001; 
      13'd2182: data <=16'b0000000001000011; 
      13'd2183: data <=16'b1111111111100111; 
      13'd2184: data <=16'b0000000000011011; 
      13'd2185: data <=16'b1111111110101010; 
      13'd2186: data <=16'b1111111100100010; 
      13'd2187: data <=16'b0000000011000011; 
      13'd2188: data <=16'b1111111110101101; 
      13'd2189: data <=16'b0000000000000100; 
      13'd2190: data <=16'b1111111101110101; 
      13'd2191: data <=16'b1111111111100011; 
      13'd2192: data <=16'b0000000000001010; 
      13'd2193: data <=16'b0000000001010000; 
      13'd2194: data <=16'b1111111110100001; 
      13'd2195: data <=16'b1111111111100110; 
      13'd2196: data <=16'b0000000000111110; 
      13'd2197: data <=16'b1111111110011100; 
      13'd2198: data <=16'b0000000001001011; 
      13'd2199: data <=16'b0000000000111110; 
      13'd2200: data <=16'b0000000001001001; 
      13'd2201: data <=16'b0000000001000010; 
      13'd2202: data <=16'b1111111110110010; 
      13'd2203: data <=16'b1111111110110010; 
      13'd2204: data <=16'b1111111111111100; 
      13'd2205: data <=16'b1111111101010101; 
      13'd2206: data <=16'b0000000000110111; 
      13'd2207: data <=16'b0000000000000110; 
      13'd2208: data <=16'b1111111111010001; 
      13'd2209: data <=16'b1111111111001100; 
      13'd2210: data <=16'b1111111110000011; 
      13'd2211: data <=16'b1111111110110110; 
      13'd2212: data <=16'b0000000000100011; 
      13'd2213: data <=16'b0000000001100111; 
      13'd2214: data <=16'b0000000001100010; 
      13'd2215: data <=16'b1111111110001110; 
      13'd2216: data <=16'b0000000000000100; 
      13'd2217: data <=16'b1111111101110001; 
      13'd2218: data <=16'b0000000000110000; 
      13'd2219: data <=16'b1111111110101000; 
      13'd2220: data <=16'b1111111100101101; 
      13'd2221: data <=16'b0000000010010110; 
      13'd2222: data <=16'b1111111110101010; 
      13'd2223: data <=16'b0000000001110111; 
      13'd2224: data <=16'b1111111110010111; 
      13'd2225: data <=16'b0000000001010101; 
      13'd2226: data <=16'b1111111111111001; 
      13'd2227: data <=16'b1111111111111000; 
      13'd2228: data <=16'b1111111111111110; 
      13'd2229: data <=16'b0000000001100110; 
      13'd2230: data <=16'b0000000010011011; 
      13'd2231: data <=16'b0000000001110001; 
      13'd2232: data <=16'b1111111111111111; 
      13'd2233: data <=16'b1111111110100110; 
      13'd2234: data <=16'b1111111111111011; 
      13'd2235: data <=16'b0000000000000010; 
      13'd2236: data <=16'b1111111111101111; 
      13'd2237: data <=16'b1111111111110011; 
      13'd2238: data <=16'b1111111110001011; 
      13'd2239: data <=16'b0000000001100110; 
      13'd2240: data <=16'b1111111111111001; 
      13'd2241: data <=16'b0000000001100010; 
      13'd2242: data <=16'b0000000000011110; 
      13'd2243: data <=16'b1111111111111100; 
      13'd2244: data <=16'b0000000001011011; 
      13'd2245: data <=16'b1111111110110110; 
      13'd2246: data <=16'b1111111111101001; 
      13'd2247: data <=16'b1111111111001001; 
      13'd2248: data <=16'b0000000010110000; 
      13'd2249: data <=16'b1111111110001011; 
      13'd2250: data <=16'b0000000010111100; 
      13'd2251: data <=16'b0000000000100010; 
      13'd2252: data <=16'b0000000000000000; 
      13'd2253: data <=16'b0000000001100010; 
      13'd2254: data <=16'b1111111111100101; 
      13'd2255: data <=16'b0000000001011111; 
      13'd2256: data <=16'b0000000000011101; 
      13'd2257: data <=16'b1111111110101110; 
      13'd2258: data <=16'b0000000000111010; 
      13'd2259: data <=16'b0000000000101100; 
      13'd2260: data <=16'b0000000010100101; 
      13'd2261: data <=16'b1111111111110101; 
      13'd2262: data <=16'b0000000000110011; 
      13'd2263: data <=16'b1111111111101011; 
      13'd2264: data <=16'b0000000000101100; 
      13'd2265: data <=16'b1111111111011100; 
      13'd2266: data <=16'b1111111100111101; 
      13'd2267: data <=16'b0000000001000000; 
      13'd2268: data <=16'b0000000001001000; 
      13'd2269: data <=16'b0000000000110101; 
      13'd2270: data <=16'b0000000010000111; 
      13'd2271: data <=16'b0000000001110001; 
      13'd2272: data <=16'b1111111111010100; 
      13'd2273: data <=16'b0000000010100011; 
      13'd2274: data <=16'b1111111111010100; 
      13'd2275: data <=16'b0000000001001010; 
      13'd2276: data <=16'b1111111100100111; 
      13'd2277: data <=16'b1111111111010010; 
      13'd2278: data <=16'b0000000001000010; 
      13'd2279: data <=16'b1111111101101101; 
      13'd2280: data <=16'b0000000000000111; 
      13'd2281: data <=16'b1111111111110001; 
      13'd2282: data <=16'b1111111101110001; 
      13'd2283: data <=16'b1111111111110100; 
      13'd2284: data <=16'b0000000000001010; 
      13'd2285: data <=16'b0000000000000101; 
      13'd2286: data <=16'b1111111110110011; 
      13'd2287: data <=16'b0000000010010100; 
      13'd2288: data <=16'b1111111111110110; 
      13'd2289: data <=16'b0000000001111101; 
      13'd2290: data <=16'b1111111111010101; 
      13'd2291: data <=16'b0000000000111010; 
      13'd2292: data <=16'b0000000000110001; 
      13'd2293: data <=16'b0000000000110110; 
      13'd2294: data <=16'b1111111111110001; 
      13'd2295: data <=16'b1111111111000001; 
      13'd2296: data <=16'b1111111101101010; 
      13'd2297: data <=16'b1111111111100000; 
      13'd2298: data <=16'b0000000000100000; 
      13'd2299: data <=16'b1111111111101011; 
      13'd2300: data <=16'b1111111110110001; 
      13'd2301: data <=16'b0000000000001011; 
      13'd2302: data <=16'b1111111110000000; 
      13'd2303: data <=16'b1111111110111111; 
      13'd2304: data <=16'b0000000001001010; 
      13'd2305: data <=16'b0000000000000110; 
      13'd2306: data <=16'b0000000001111011; 
      13'd2307: data <=16'b0000000010011001; 
      13'd2308: data <=16'b0000000010001000; 
      13'd2309: data <=16'b1111111100001101; 
      13'd2310: data <=16'b1111111110100010; 
      13'd2311: data <=16'b1111111110100100; 
      13'd2312: data <=16'b0000000000110111; 
      13'd2313: data <=16'b0000000000100100; 
      13'd2314: data <=16'b0000000000010010; 
      13'd2315: data <=16'b0000000000101010; 
      13'd2316: data <=16'b0000000000101001; 
      13'd2317: data <=16'b1111111110100111; 
      13'd2318: data <=16'b0000000000110111; 
      13'd2319: data <=16'b0000000001110100; 
      13'd2320: data <=16'b1111111111001110; 
      13'd2321: data <=16'b0000000001111101; 
      13'd2322: data <=16'b0000000001011010; 
      13'd2323: data <=16'b1111111101011011; 
      13'd2324: data <=16'b1111111111011100; 
      13'd2325: data <=16'b1111111110000011; 
      13'd2326: data <=16'b0000000000100111; 
      13'd2327: data <=16'b0000000000111001; 
      13'd2328: data <=16'b1111111100110110; 
      13'd2329: data <=16'b0000000001000100; 
      13'd2330: data <=16'b1111111111110010; 
      13'd2331: data <=16'b0000000000000011; 
      13'd2332: data <=16'b1111111111101001; 
      13'd2333: data <=16'b1111111110001010; 
      13'd2334: data <=16'b0000000000101011; 
      13'd2335: data <=16'b0000000001000110; 
      13'd2336: data <=16'b0000000010110010; 
      13'd2337: data <=16'b1111111111101010; 
      13'd2338: data <=16'b1111111111101100; 
      13'd2339: data <=16'b1111111101110110; 
      13'd2340: data <=16'b1111111110111111; 
      13'd2341: data <=16'b1111111110101110; 
      13'd2342: data <=16'b1111111111111111; 
      13'd2343: data <=16'b0000000001001110; 
      13'd2344: data <=16'b1111111111000011; 
      13'd2345: data <=16'b1111111110001100; 
      13'd2346: data <=16'b0000000010100101; 
      13'd2347: data <=16'b0000000001111011; 
      13'd2348: data <=16'b1111111111001111; 
      13'd2349: data <=16'b1111111111010010; 
      13'd2350: data <=16'b0000000000011011; 
      13'd2351: data <=16'b1111111110111001; 
      13'd2352: data <=16'b1111111111001100; 
      13'd2353: data <=16'b0000000000011110; 
      13'd2354: data <=16'b1111111111100110; 
      13'd2355: data <=16'b0000000001000101; 
      13'd2356: data <=16'b0000000010011010; 
      13'd2357: data <=16'b1111111110111010; 
      13'd2358: data <=16'b1111111110100111; 
      13'd2359: data <=16'b1111111110110011; 
      13'd2360: data <=16'b1111111111110111; 
      13'd2361: data <=16'b1111111101101101; 
      13'd2362: data <=16'b1111111111011110; 
      13'd2363: data <=16'b1111111100111100; 
      13'd2364: data <=16'b0000000000010000; 
      13'd2365: data <=16'b0000000000111010; 
      13'd2366: data <=16'b1111111101000101; 
      13'd2367: data <=16'b1111111111111001; 
      13'd2368: data <=16'b1111111111100000; 
      13'd2369: data <=16'b0000000010010101; 
      13'd2370: data <=16'b1111111111010111; 
      13'd2371: data <=16'b0000000000010010; 
      13'd2372: data <=16'b1111111111111101; 
      13'd2373: data <=16'b1111111111010011; 
      13'd2374: data <=16'b1111111101111001; 
      13'd2375: data <=16'b0000000001101011; 
      13'd2376: data <=16'b0000000000001001; 
      13'd2377: data <=16'b0000000001000100; 
      13'd2378: data <=16'b0000000001111001; 
      13'd2379: data <=16'b0000000001001001; 
      13'd2380: data <=16'b0000000010001111; 
      13'd2381: data <=16'b1111111110001010; 
      13'd2382: data <=16'b0000000000000001; 
      13'd2383: data <=16'b1111111110110110; 
      13'd2384: data <=16'b1111111101011110; 
      13'd2385: data <=16'b1111111111001010; 
      13'd2386: data <=16'b0000000000010101; 
      13'd2387: data <=16'b0000000000011000; 
      13'd2388: data <=16'b1111111111000000; 
      13'd2389: data <=16'b0000000000001110; 
      13'd2390: data <=16'b0000000010010111; 
      13'd2391: data <=16'b1111111110001001; 
      13'd2392: data <=16'b1111111110110000; 
      13'd2393: data <=16'b0000000000101011; 
      13'd2394: data <=16'b0000000010000100; 
      13'd2395: data <=16'b1111111111101001; 
      13'd2396: data <=16'b0000000010111110; 
      13'd2397: data <=16'b0000000001000110; 
      13'd2398: data <=16'b1111111111011011; 
      13'd2399: data <=16'b0000000001010000; 
      13'd2400: data <=16'b0000000000000100; 
      13'd2401: data <=16'b1111111111000110; 
      13'd2402: data <=16'b0000000000000101; 
      13'd2403: data <=16'b0000000001011010; 
      13'd2404: data <=16'b0000000001011011; 
      13'd2405: data <=16'b1111111111011011; 
      13'd2406: data <=16'b1111111110110110; 
      13'd2407: data <=16'b1111111110110111; 
      13'd2408: data <=16'b0000000000000111; 
      13'd2409: data <=16'b0000000000000011; 
      13'd2410: data <=16'b0000000010110000; 
      13'd2411: data <=16'b0000000000011100; 
      13'd2412: data <=16'b1111111111001100; 
      13'd2413: data <=16'b0000000001111011; 
      13'd2414: data <=16'b0000000000101100; 
      13'd2415: data <=16'b0000000001100001; 
      13'd2416: data <=16'b1111111110011010; 
      13'd2417: data <=16'b0000000010110010; 
      13'd2418: data <=16'b1111111101011100; 
      13'd2419: data <=16'b0000000010010111; 
      13'd2420: data <=16'b1111111110001001; 
      13'd2421: data <=16'b1111111111100010; 
      13'd2422: data <=16'b0000000000100000; 
      13'd2423: data <=16'b1111111111110110; 
      13'd2424: data <=16'b1111111111111110; 
      13'd2425: data <=16'b0000000000100011; 
      13'd2426: data <=16'b1111111101110000; 
      13'd2427: data <=16'b1111111110110100; 
      13'd2428: data <=16'b1111111111110100; 
      13'd2429: data <=16'b0000000000010001; 
      13'd2430: data <=16'b1111111111111100; 
      13'd2431: data <=16'b1111111110100010; 
      13'd2432: data <=16'b0000000000101101; 
      13'd2433: data <=16'b0000000000000011; 
      13'd2434: data <=16'b1111111111101100; 
      13'd2435: data <=16'b0000000001000100; 
      13'd2436: data <=16'b1111111110001010; 
      13'd2437: data <=16'b0000000001111111; 
      13'd2438: data <=16'b1111111111001111; 
      13'd2439: data <=16'b0000000001010111; 
      13'd2440: data <=16'b1111111111010000; 
      13'd2441: data <=16'b0000000000111001; 
      13'd2442: data <=16'b1111111101100111; 
      13'd2443: data <=16'b0000000000111100; 
      13'd2444: data <=16'b0000000010110011; 
      13'd2445: data <=16'b0000000000010101; 
      13'd2446: data <=16'b1111111111011110; 
      13'd2447: data <=16'b0000000000110100; 
      13'd2448: data <=16'b1111111110100111; 
      13'd2449: data <=16'b1111111110100100; 
      13'd2450: data <=16'b0000000000010001; 
      13'd2451: data <=16'b1111111111110110; 
      13'd2452: data <=16'b1111111111100111; 
      13'd2453: data <=16'b0000000001001000; 
      13'd2454: data <=16'b1111111111001001; 
      13'd2455: data <=16'b0000000000011100; 
      13'd2456: data <=16'b1111111111100111; 
      13'd2457: data <=16'b0000000001011011; 
      13'd2458: data <=16'b1111111111001011; 
      13'd2459: data <=16'b1111111101100101; 
      13'd2460: data <=16'b1111111111100111; 
      13'd2461: data <=16'b0000000001011010; 
      13'd2462: data <=16'b1111111111000001; 
      13'd2463: data <=16'b1111111110111000; 
      13'd2464: data <=16'b1111111111011100; 
      13'd2465: data <=16'b1111111110110110; 
      13'd2466: data <=16'b1111111111001010; 
      13'd2467: data <=16'b0000000010010100; 
      13'd2468: data <=16'b1111111110111100; 
      13'd2469: data <=16'b1111111110011000; 
      13'd2470: data <=16'b0000000000101011; 
      13'd2471: data <=16'b1111111101101101; 
      13'd2472: data <=16'b0000000001100001; 
      13'd2473: data <=16'b0000000000011010; 
      13'd2474: data <=16'b1111111111111011; 
      13'd2475: data <=16'b0000000000110001; 
      13'd2476: data <=16'b0000000001000000; 
      13'd2477: data <=16'b0000000000010000; 
      13'd2478: data <=16'b0000000001100110; 
      13'd2479: data <=16'b1111111111011100; 
      13'd2480: data <=16'b1111111101101111; 
      13'd2481: data <=16'b0000000000011101; 
      13'd2482: data <=16'b0000000001110110; 
      13'd2483: data <=16'b1111111110010001; 
      13'd2484: data <=16'b1111111110000011; 
      13'd2485: data <=16'b1111111111110111; 
      13'd2486: data <=16'b0000000001001000; 
      13'd2487: data <=16'b0000000010000000; 
      13'd2488: data <=16'b1111111110001111; 
      13'd2489: data <=16'b1111111111111110; 
      13'd2490: data <=16'b0000000001101001; 
      13'd2491: data <=16'b0000000000101100; 
      13'd2492: data <=16'b1111111110010011; 
      13'd2493: data <=16'b0000000001000111; 
      13'd2494: data <=16'b1111111111011010; 
      13'd2495: data <=16'b0000000001000001; 
      13'd2496: data <=16'b0000000000101110; 
      13'd2497: data <=16'b0000000000001001; 
      13'd2498: data <=16'b1111111111001010; 
      13'd2499: data <=16'b1111111110011100; 
      13'd2500: data <=16'b0000000010001110; 
      13'd2501: data <=16'b1111111111001100; 
      13'd2502: data <=16'b0000000011001011; 
      13'd2503: data <=16'b0000000000100100; 
      13'd2504: data <=16'b0000000000101000; 
      13'd2505: data <=16'b0000000001110110; 
      13'd2506: data <=16'b0000000000100101; 
      13'd2507: data <=16'b1111111110111000; 
      13'd2508: data <=16'b0000000000001001; 
      13'd2509: data <=16'b1111111111101111; 
      13'd2510: data <=16'b1111111101101111; 
      13'd2511: data <=16'b0000000000101011; 
      13'd2512: data <=16'b0000000000100101; 
      13'd2513: data <=16'b0000000000011110; 
      13'd2514: data <=16'b1111111101001101; 
      13'd2515: data <=16'b0000000001110010; 
      13'd2516: data <=16'b0000000000101000; 
      13'd2517: data <=16'b0000000010001110; 
      13'd2518: data <=16'b0000000000010011; 
      13'd2519: data <=16'b1111111111001010; 
      13'd2520: data <=16'b0000000000000000; 
      13'd2521: data <=16'b0000000000000001; 
      13'd2522: data <=16'b0000000001101010; 
      13'd2523: data <=16'b0000000001111101; 
      13'd2524: data <=16'b1111111111000001; 
      13'd2525: data <=16'b0000000000001100; 
      13'd2526: data <=16'b0000000000000001; 
      13'd2527: data <=16'b1111111111110100; 
      13'd2528: data <=16'b1111111110101011; 
      13'd2529: data <=16'b0000000011101111; 
      13'd2530: data <=16'b1111111111101000; 
      13'd2531: data <=16'b0000000010011100; 
      13'd2532: data <=16'b1111111110110100; 
      13'd2533: data <=16'b0000000000101100; 
      13'd2534: data <=16'b0000000000011000; 
      13'd2535: data <=16'b0000000010110000; 
      13'd2536: data <=16'b0000000000000001; 
      13'd2537: data <=16'b1111111111100111; 
      13'd2538: data <=16'b1111111101000100; 
      13'd2539: data <=16'b0000000000010100; 
      13'd2540: data <=16'b1111111011110101; 
      13'd2541: data <=16'b0000000000000000; 
      13'd2542: data <=16'b0000000000111011; 
      13'd2543: data <=16'b0000000000111100; 
      13'd2544: data <=16'b1111111110011110; 
      13'd2545: data <=16'b0000000001010011; 
      13'd2546: data <=16'b0000000001101011; 
      13'd2547: data <=16'b0000000010001101; 
      13'd2548: data <=16'b0000000000110100; 
      13'd2549: data <=16'b1111111111101000; 
      13'd2550: data <=16'b0000000000011101; 
      13'd2551: data <=16'b1111111110111111; 
      13'd2552: data <=16'b1111111111101110; 
      13'd2553: data <=16'b1111111110011101; 
      13'd2554: data <=16'b0000000000011101; 
      13'd2555: data <=16'b1111111111001100; 
      13'd2556: data <=16'b1111111110111000; 
      13'd2557: data <=16'b0000000000010010; 
      13'd2558: data <=16'b1111111101000011; 
      13'd2559: data <=16'b0000000000011110; 
      13'd2560: data <=16'b0000000000110001; 
      13'd2561: data <=16'b0000000000001010; 
      13'd2562: data <=16'b0000000000011101; 
      13'd2563: data <=16'b0000000000111001; 
      13'd2564: data <=16'b1111111101111111; 
      13'd2565: data <=16'b1111111111011100; 
      13'd2566: data <=16'b1111111111110111; 
      13'd2567: data <=16'b1111111110001101; 
      13'd2568: data <=16'b0000000001000011; 
      13'd2569: data <=16'b1111111110011100; 
      13'd2570: data <=16'b1111111110110011; 
      13'd2571: data <=16'b0000000000001100; 
      13'd2572: data <=16'b1111111111010111; 
      13'd2573: data <=16'b0000000000010111; 
      13'd2574: data <=16'b1111111111000001; 
      13'd2575: data <=16'b0000000010110100; 
      13'd2576: data <=16'b0000000001101011; 
      13'd2577: data <=16'b0000000001100110; 
      13'd2578: data <=16'b1111111101000111; 
      13'd2579: data <=16'b1111111110110111; 
      13'd2580: data <=16'b1111111111000110; 
      13'd2581: data <=16'b1111111111001011; 
      13'd2582: data <=16'b1111111111011001; 
      13'd2583: data <=16'b0000000000010111; 
      13'd2584: data <=16'b1111111111011110; 
      13'd2585: data <=16'b0000000000110010; 
      13'd2586: data <=16'b1111111111001001; 
      13'd2587: data <=16'b1111111100111101; 
      13'd2588: data <=16'b0000000000000010; 
      13'd2589: data <=16'b0000000000001010; 
      13'd2590: data <=16'b0000000000010001; 
      13'd2591: data <=16'b0000000001001111; 
      13'd2592: data <=16'b0000000000001101; 
      13'd2593: data <=16'b1111111101000001; 
      13'd2594: data <=16'b1111111110111011; 
      13'd2595: data <=16'b0000000000001001; 
      13'd2596: data <=16'b0000000010000101; 
      13'd2597: data <=16'b1111111111111110; 
      13'd2598: data <=16'b1111111111001011; 
      13'd2599: data <=16'b0000000010011101; 
      13'd2600: data <=16'b1111111111000101; 
      13'd2601: data <=16'b0000000000011010; 
      13'd2602: data <=16'b1111111110101001; 
      13'd2603: data <=16'b0000000000111010; 
      13'd2604: data <=16'b0000000010010000; 
      13'd2605: data <=16'b1111111111111010; 
      13'd2606: data <=16'b1111111110110011; 
      13'd2607: data <=16'b1111111101011000; 
      13'd2608: data <=16'b1111111111101101; 
      13'd2609: data <=16'b1111111110100001; 
      13'd2610: data <=16'b1111111111111000; 
      13'd2611: data <=16'b1111111100101101; 
      13'd2612: data <=16'b1111111111101011; 
      13'd2613: data <=16'b1111111110110111; 
      13'd2614: data <=16'b1111111111111001; 
      13'd2615: data <=16'b1111111111011011; 
      13'd2616: data <=16'b1111111110100110; 
      13'd2617: data <=16'b0000000000100111; 
      13'd2618: data <=16'b0000000000001101; 
      13'd2619: data <=16'b0000000000010010; 
      13'd2620: data <=16'b1111111111001000; 
      13'd2621: data <=16'b1111111101100101; 
      13'd2622: data <=16'b1111111111000101; 
      13'd2623: data <=16'b0000000001101110; 
      13'd2624: data <=16'b0000000000001001; 
      13'd2625: data <=16'b0000000001100100; 
      13'd2626: data <=16'b1111111111001111; 
      13'd2627: data <=16'b1111111111101000; 
      13'd2628: data <=16'b0000000000101110; 
      13'd2629: data <=16'b1111111100110111; 
      13'd2630: data <=16'b1111111101100010; 
      13'd2631: data <=16'b1111111111100101; 
      13'd2632: data <=16'b1111111111011010; 
      13'd2633: data <=16'b0000000010010001; 
      13'd2634: data <=16'b0000000000110110; 
      13'd2635: data <=16'b1111111101111001; 
      13'd2636: data <=16'b0000000000100101; 
      13'd2637: data <=16'b0000000001010110; 
      13'd2638: data <=16'b0000000000100100; 
      13'd2639: data <=16'b0000000000100101; 
      13'd2640: data <=16'b0000000000011011; 
      13'd2641: data <=16'b1111111101001001; 
      13'd2642: data <=16'b0000000000000010; 
      13'd2643: data <=16'b0000000000101010; 
      13'd2644: data <=16'b1111111110011010; 
      13'd2645: data <=16'b0000000000010101; 
      13'd2646: data <=16'b1111111111101111; 
      13'd2647: data <=16'b0000000001011011; 
      13'd2648: data <=16'b1111111110100011; 
      13'd2649: data <=16'b1111111101011110; 
      13'd2650: data <=16'b0000000001001111; 
      13'd2651: data <=16'b1111111111100010; 
      13'd2652: data <=16'b1111111111111100; 
      13'd2653: data <=16'b1111111110111011; 
      13'd2654: data <=16'b0000000000111001; 
      13'd2655: data <=16'b1111111111101111; 
      13'd2656: data <=16'b0000000001011011; 
      13'd2657: data <=16'b1111111111111001; 
      13'd2658: data <=16'b1111111111100011; 
      13'd2659: data <=16'b1111111111111000; 
      13'd2660: data <=16'b0000000001100011; 
      13'd2661: data <=16'b0000000001001111; 
      13'd2662: data <=16'b1111111101110000; 
      13'd2663: data <=16'b0000000000111101; 
      13'd2664: data <=16'b1111111011001110; 
      13'd2665: data <=16'b0000000000110001; 
      13'd2666: data <=16'b1111111110100100; 
      13'd2667: data <=16'b0000000001010011; 
      13'd2668: data <=16'b1111111101101010; 
      13'd2669: data <=16'b1111111111010000; 
      13'd2670: data <=16'b1111111110101010; 
      13'd2671: data <=16'b0000000000001110; 
      13'd2672: data <=16'b0000000001010011; 
      13'd2673: data <=16'b0000000010001100; 
      13'd2674: data <=16'b0000000001000101; 
      13'd2675: data <=16'b1111111110101011; 
      13'd2676: data <=16'b0000000000101010; 
      13'd2677: data <=16'b0000000000011011; 
      13'd2678: data <=16'b0000000011100100; 
      13'd2679: data <=16'b0000000000010111; 
      13'd2680: data <=16'b1111111111010011; 
      13'd2681: data <=16'b1111111111000010; 
      13'd2682: data <=16'b0000000000000100; 
      13'd2683: data <=16'b0000000001110100; 
      13'd2684: data <=16'b0000000000001010; 
      13'd2685: data <=16'b1111111111101100; 
      13'd2686: data <=16'b0000000000000000; 
      13'd2687: data <=16'b1111111101011100; 
      13'd2688: data <=16'b1111111111111100; 
      13'd2689: data <=16'b0000000000111111; 
      13'd2690: data <=16'b0000000001000001; 
      13'd2691: data <=16'b1111111111011101; 
      13'd2692: data <=16'b1111111101111100; 
      13'd2693: data <=16'b1111111111001100; 
      13'd2694: data <=16'b1111111110100011; 
      13'd2695: data <=16'b1111111110011101; 
      13'd2696: data <=16'b0000000010000000; 
      13'd2697: data <=16'b0000000000101100; 
      13'd2698: data <=16'b1111111110011110; 
      13'd2699: data <=16'b1111111111110110; 
      13'd2700: data <=16'b1111111110011110; 
      13'd2701: data <=16'b0000000011001111; 
      13'd2702: data <=16'b1111111110011000; 
      13'd2703: data <=16'b0000000001001000; 
      13'd2704: data <=16'b0000000000000110; 
      13'd2705: data <=16'b1111111110001010; 
      13'd2706: data <=16'b0000000001000111; 
      13'd2707: data <=16'b0000000100111111; 
      13'd2708: data <=16'b0000000010100111; 
      13'd2709: data <=16'b1111111111111011; 
      13'd2710: data <=16'b0000000010000000; 
      13'd2711: data <=16'b1111111111100110; 
      13'd2712: data <=16'b1111111110101001; 
      13'd2713: data <=16'b0000000000101011; 
      13'd2714: data <=16'b0000000000001010; 
      13'd2715: data <=16'b0000000000000110; 
      13'd2716: data <=16'b0000000000011100; 
      13'd2717: data <=16'b0000000010111101; 
      13'd2718: data <=16'b1111111111111011; 
      13'd2719: data <=16'b1111111111101001; 
      13'd2720: data <=16'b0000000000010111; 
      13'd2721: data <=16'b0000000000111001; 
      13'd2722: data <=16'b0000000001110011; 
      13'd2723: data <=16'b0000000000111011; 
      13'd2724: data <=16'b0000000000000001; 
      13'd2725: data <=16'b0000000000101011; 
      13'd2726: data <=16'b0000000001000110; 
      13'd2727: data <=16'b1111111111110011; 
      13'd2728: data <=16'b1111111111110101; 
      13'd2729: data <=16'b1111111111100010; 
      13'd2730: data <=16'b0000000001001010; 
      13'd2731: data <=16'b0000000010000110; 
      13'd2732: data <=16'b0000000001100110; 
      13'd2733: data <=16'b1111111111001011; 
      13'd2734: data <=16'b1111111111100010; 
      13'd2735: data <=16'b0000000001011001; 
      13'd2736: data <=16'b1111111111000110; 
      13'd2737: data <=16'b0000000001101010; 
      13'd2738: data <=16'b1111111111001010; 
      13'd2739: data <=16'b0000000000101011; 
      13'd2740: data <=16'b1111111110101001; 
      13'd2741: data <=16'b1111111101111001; 
      13'd2742: data <=16'b0000000000111100; 
      13'd2743: data <=16'b0000000011111000; 
      13'd2744: data <=16'b0000000001000000; 
      13'd2745: data <=16'b1111111111110001; 
      13'd2746: data <=16'b0000000011011000; 
      13'd2747: data <=16'b1111111101111011; 
      13'd2748: data <=16'b0000000000011110; 
      13'd2749: data <=16'b1111111111010101; 
      13'd2750: data <=16'b0000000010110010; 
      13'd2751: data <=16'b0000000010001010; 
      13'd2752: data <=16'b0000000001001110; 
      13'd2753: data <=16'b0000000001110101; 
      13'd2754: data <=16'b0000000010010000; 
      13'd2755: data <=16'b1111111101110001; 
      13'd2756: data <=16'b0000000010000110; 
      13'd2757: data <=16'b1111111111101011; 
      13'd2758: data <=16'b0000000001111001; 
      13'd2759: data <=16'b0000000000001111; 
      13'd2760: data <=16'b0000000001001001; 
      13'd2761: data <=16'b0000000010010111; 
      13'd2762: data <=16'b1111111111000001; 
      13'd2763: data <=16'b0000000000111010; 
      13'd2764: data <=16'b0000000000011100; 
      13'd2765: data <=16'b0000000000010010; 
      13'd2766: data <=16'b1111111111111101; 
      13'd2767: data <=16'b0000000001100001; 
      13'd2768: data <=16'b0000000000101011; 
      13'd2769: data <=16'b1111111110010001; 
      13'd2770: data <=16'b0000000001000000; 
      13'd2771: data <=16'b1111111111100111; 
      13'd2772: data <=16'b0000000001111010; 
      13'd2773: data <=16'b0000000010000110; 
      13'd2774: data <=16'b0000000010110000; 
      13'd2775: data <=16'b1111111110110001; 
      13'd2776: data <=16'b0000000000110110; 
      13'd2777: data <=16'b1111111101111101; 
      13'd2778: data <=16'b0000000011000100; 
      13'd2779: data <=16'b1111111111101110; 
      13'd2780: data <=16'b1111111111001101; 
      13'd2781: data <=16'b0000000000001011; 
      13'd2782: data <=16'b0000000010100010; 
      13'd2783: data <=16'b0000000000010010; 
      13'd2784: data <=16'b0000000001011010; 
      13'd2785: data <=16'b1111111111001111; 
      13'd2786: data <=16'b0000000001001001; 
      13'd2787: data <=16'b0000000010101100; 
      13'd2788: data <=16'b0000000001000001; 
      13'd2789: data <=16'b0000000000000111; 
      13'd2790: data <=16'b0000000000100010; 
      13'd2791: data <=16'b0000000000001001; 
      13'd2792: data <=16'b1111111101101011; 
      13'd2793: data <=16'b1111111111000011; 
      13'd2794: data <=16'b0000000001001010; 
      13'd2795: data <=16'b1111111101010110; 
      13'd2796: data <=16'b1111111101001111; 
      13'd2797: data <=16'b1111111111000010; 
      13'd2798: data <=16'b1111111111110000; 
      13'd2799: data <=16'b1111111101001011; 
      13'd2800: data <=16'b1111111111100010; 
      13'd2801: data <=16'b1111111110110111; 
      13'd2802: data <=16'b0000000000101110; 
      13'd2803: data <=16'b0000000100010000; 
      13'd2804: data <=16'b0000000000101010; 
      13'd2805: data <=16'b1111111110111100; 
      13'd2806: data <=16'b0000000000001110; 
      13'd2807: data <=16'b1111111111010100; 
      13'd2808: data <=16'b0000000000001111; 
      13'd2809: data <=16'b1111111110100101; 
      13'd2810: data <=16'b0000000001110010; 
      13'd2811: data <=16'b0000000001011010; 
      13'd2812: data <=16'b0000000001100111; 
      13'd2813: data <=16'b0000000001100000; 
      13'd2814: data <=16'b0000000001000001; 
      13'd2815: data <=16'b0000000010010100; 
      13'd2816: data <=16'b0000000000111010; 
      13'd2817: data <=16'b0000000001101110; 
      13'd2818: data <=16'b1111111111111111; 
      13'd2819: data <=16'b0000000010111111; 
      13'd2820: data <=16'b0000000000011000; 
      13'd2821: data <=16'b1111111110100101; 
      13'd2822: data <=16'b1111111111001100; 
      13'd2823: data <=16'b1111111111110000; 
      13'd2824: data <=16'b0000000001111010; 
      13'd2825: data <=16'b1111111111000110; 
      13'd2826: data <=16'b1111111111100101; 
      13'd2827: data <=16'b1111111111011100; 
      13'd2828: data <=16'b1111111111001110; 
      13'd2829: data <=16'b0000000001100111; 
      13'd2830: data <=16'b1111111101111011; 
      13'd2831: data <=16'b1111111110100000; 
      13'd2832: data <=16'b1111111110011001; 
      13'd2833: data <=16'b0000000000101101; 
      13'd2834: data <=16'b1111111101110010; 
      13'd2835: data <=16'b0000000000111000; 
      13'd2836: data <=16'b0000000000100100; 
      13'd2837: data <=16'b1111111111010011; 
      13'd2838: data <=16'b0000000000011110; 
      13'd2839: data <=16'b0000000001001000; 
      13'd2840: data <=16'b1111111111100110; 
      13'd2841: data <=16'b1111111111011101; 
      13'd2842: data <=16'b0000000000001001; 
      13'd2843: data <=16'b1111111110100110; 
      13'd2844: data <=16'b1111111110101101; 
      13'd2845: data <=16'b1111111111001100; 
      13'd2846: data <=16'b0000000001000010; 
      13'd2847: data <=16'b1111111111101101; 
      13'd2848: data <=16'b0000000000010001; 
      13'd2849: data <=16'b1111111101110101; 
      13'd2850: data <=16'b1111111110100000; 
      13'd2851: data <=16'b1111111111100001; 
      13'd2852: data <=16'b1111111110100101; 
      13'd2853: data <=16'b1111111110110101; 
      13'd2854: data <=16'b1111111110110100; 
      13'd2855: data <=16'b0000000011001000; 
      13'd2856: data <=16'b0000000010101100; 
      13'd2857: data <=16'b0000000000000001; 
      13'd2858: data <=16'b0000000010001110; 
      13'd2859: data <=16'b0000000001100000; 
      13'd2860: data <=16'b1111111111111001; 
      13'd2861: data <=16'b0000000000000001; 
      13'd2862: data <=16'b0000000000001101; 
      13'd2863: data <=16'b1111111111111001; 
      13'd2864: data <=16'b0000000001011011; 
      13'd2865: data <=16'b1111111110101100; 
      13'd2866: data <=16'b1111111111101001; 
      13'd2867: data <=16'b1111111111010101; 
      13'd2868: data <=16'b0000000001100111; 
      13'd2869: data <=16'b1111111110101101; 
      13'd2870: data <=16'b1111111110101011; 
      13'd2871: data <=16'b0000000000101110; 
      13'd2872: data <=16'b1111111110001001; 
      13'd2873: data <=16'b1111111110110011; 
      13'd2874: data <=16'b0000000001100100; 
      13'd2875: data <=16'b0000000000110010; 
      13'd2876: data <=16'b0000000001001111; 
      13'd2877: data <=16'b1111111110111010; 
      13'd2878: data <=16'b1111111111101000; 
      13'd2879: data <=16'b0000000000011110; 
      13'd2880: data <=16'b1111111101101111; 
      13'd2881: data <=16'b0000000000101100; 
      13'd2882: data <=16'b1111111110100110; 
      13'd2883: data <=16'b0000000001001100; 
      13'd2884: data <=16'b0000000000110001; 
      13'd2885: data <=16'b1111111111001100; 
      13'd2886: data <=16'b0000000000101011; 
      13'd2887: data <=16'b1111111111000000; 
      13'd2888: data <=16'b1111111110001111; 
      13'd2889: data <=16'b1111111110110101; 
      13'd2890: data <=16'b0000000001011000; 
      13'd2891: data <=16'b0000000001011110; 
      13'd2892: data <=16'b1111111111101101; 
      13'd2893: data <=16'b0000000000101110; 
      13'd2894: data <=16'b1111111100010110; 
      13'd2895: data <=16'b1111111111010001; 
      13'd2896: data <=16'b1111111111101111; 
      13'd2897: data <=16'b0000000000101111; 
      13'd2898: data <=16'b0000000000110010; 
      13'd2899: data <=16'b0000000000100111; 
      13'd2900: data <=16'b1111111111001000; 
      13'd2901: data <=16'b1111111111100111; 
      13'd2902: data <=16'b0000000001010110; 
      13'd2903: data <=16'b1111111101111010; 
      13'd2904: data <=16'b0000000000111110; 
      13'd2905: data <=16'b0000000000000010; 
      13'd2906: data <=16'b0000000000100011; 
      13'd2907: data <=16'b0000000010000001; 
      13'd2908: data <=16'b1111111111000111; 
      13'd2909: data <=16'b1111111110001010; 
      13'd2910: data <=16'b1111111111001100; 
      13'd2911: data <=16'b0000000000011000; 
      13'd2912: data <=16'b0000000010000110; 
      13'd2913: data <=16'b0000000000001011; 
      13'd2914: data <=16'b0000000001011000; 
      13'd2915: data <=16'b0000000000001000; 
      13'd2916: data <=16'b0000000000000110; 
      13'd2917: data <=16'b1111111111101011; 
      13'd2918: data <=16'b1111111100101101; 
      13'd2919: data <=16'b0000000001101110; 
      13'd2920: data <=16'b0000000001110010; 
      13'd2921: data <=16'b1111111111111011; 
      13'd2922: data <=16'b0000000000010000; 
      13'd2923: data <=16'b0000000000111001; 
      13'd2924: data <=16'b0000000000110111; 
      13'd2925: data <=16'b0000000000111110; 
      13'd2926: data <=16'b0000000000000001; 
      13'd2927: data <=16'b1111111111011110; 
      13'd2928: data <=16'b0000000001110001; 
      13'd2929: data <=16'b1111111110010100; 
      13'd2930: data <=16'b0000000010000100; 
      13'd2931: data <=16'b0000000000110110; 
      13'd2932: data <=16'b0000000001010010; 
      13'd2933: data <=16'b0000000001001111; 
      13'd2934: data <=16'b0000000011111000; 
      13'd2935: data <=16'b0000000001011010; 
      13'd2936: data <=16'b0000000001001000; 
      13'd2937: data <=16'b1111111100100010; 
      13'd2938: data <=16'b1111111110000100; 
      13'd2939: data <=16'b0000000001110011; 
      13'd2940: data <=16'b1111111111101100; 
      13'd2941: data <=16'b1111111111111111; 
      13'd2942: data <=16'b1111111111101100; 
      13'd2943: data <=16'b0000000001000111; 
      13'd2944: data <=16'b0000000000010010; 
      13'd2945: data <=16'b0000000010000101; 
      13'd2946: data <=16'b0000000010010111; 
      13'd2947: data <=16'b1111111111111000; 
      13'd2948: data <=16'b1111111101111100; 
      13'd2949: data <=16'b1111111111110010; 
      13'd2950: data <=16'b0000000001011000; 
      13'd2951: data <=16'b1111111111111000; 
      13'd2952: data <=16'b1111111110100101; 
      13'd2953: data <=16'b0000000001110101; 
      13'd2954: data <=16'b1111111110001110; 
      13'd2955: data <=16'b0000000001001001; 
      13'd2956: data <=16'b1111111101011101; 
      13'd2957: data <=16'b0000000001001011; 
      13'd2958: data <=16'b1111111101010100; 
      13'd2959: data <=16'b1111111111011111; 
      13'd2960: data <=16'b0000000000110110; 
      13'd2961: data <=16'b0000000000101111; 
      13'd2962: data <=16'b1111111110101000; 
      13'd2963: data <=16'b1111111110100000; 
      13'd2964: data <=16'b0000000000101010; 
      13'd2965: data <=16'b1111111111001001; 
      13'd2966: data <=16'b1111111111110010; 
      13'd2967: data <=16'b1111111111000011; 
      13'd2968: data <=16'b1111111110010110; 
      13'd2969: data <=16'b0000000001111001; 
      13'd2970: data <=16'b1111111110100100; 
      13'd2971: data <=16'b1111111101110011; 
      13'd2972: data <=16'b1111111111011000; 
      13'd2973: data <=16'b0000000000011011; 
      13'd2974: data <=16'b0000000001101110; 
      13'd2975: data <=16'b1111111101010000; 
      13'd2976: data <=16'b0000000001100111; 
      13'd2977: data <=16'b1111111101100011; 
      13'd2978: data <=16'b1111111111101110; 
      13'd2979: data <=16'b0000000001000000; 
      13'd2980: data <=16'b1111111101000100; 
      13'd2981: data <=16'b1111111110011000; 
      13'd2982: data <=16'b0000000001000100; 
      13'd2983: data <=16'b0000000000110010; 
      13'd2984: data <=16'b1111111111111101; 
      13'd2985: data <=16'b1111111111110010; 
      13'd2986: data <=16'b1111111101111110; 
      13'd2987: data <=16'b1111111101001011; 
      13'd2988: data <=16'b0000000011000001; 
      13'd2989: data <=16'b0000000001010011; 
      13'd2990: data <=16'b1111111111011111; 
      13'd2991: data <=16'b1111111111000010; 
      13'd2992: data <=16'b1111111111000111; 
      13'd2993: data <=16'b0000000001100011; 
      13'd2994: data <=16'b1111111111001110; 
      13'd2995: data <=16'b1111111110001110; 
      13'd2996: data <=16'b0000000000000001; 
      13'd2997: data <=16'b0000000010100000; 
      13'd2998: data <=16'b0000000000000000; 
      13'd2999: data <=16'b1111111111101011; 
      default: data<=13'd0;
    endcase 
  end 
endmodule 
